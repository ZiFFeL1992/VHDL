library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity seno_4kX20 is
port (
ADDR : std_logic_vector(11 downto 0);
CLK: std_logic;
DOUT : out std_logic_vector(19 downto 0) );
attribute rom_style         : string;
  attribute rom_style of seno_4kX20 : entity is "distributed";

end seno_4kX20;

architecture rtl of seno_4kX20 is
signal DOUT_aux : std_logic_vector(19 downto 0);
 type cell is array (0 to 4095) of std_logic_vector(19 downto 0);
constant memoria : cell :=(
0=> x"00000",
 1=> x"00324",
 2=> x"00648",
 3=> x"0096D",
 4=> x"00C91",
 5=> x"00FB6",
 6=> x"012DA",
 7=> x"015FE",
 8=> x"01923",
 9=> x"01C47",
 10=> x"01F6C",
 11=> x"02290",
 12=> x"025B4",
 13=> x"028D9",
 14=> x"02BFD",
 15=> x"02F21",
 16=> x"03245",
 17=> x"03569",
 18=> x"0388E",
 19=> x"03BB2",
 20=> x"03ED6",
 21=> x"041FA",
 22=> x"0451E",
 23=> x"04842",
 24=> x"04B66",
 25=> x"04E8A",
 26=> x"051AD",
 27=> x"054D1",
 28=> x"057F5",
 29=> x"05B19",
 30=> x"05E3C",
 31=> x"06160",
 32=> x"06483",
 33=> x"067A7",
 34=> x"06ACA",
 35=> x"06DED",
 36=> x"07111",
 37=> x"07434",
 38=> x"07757",
 39=> x"07A7A",
 40=> x"07D9D",
 41=> x"080C0",
 42=> x"083E3",
 43=> x"08705",
 44=> x"08A28",
 45=> x"08D4B",
 46=> x"0906D",
 47=> x"09390",
 48=> x"096B2",
 49=> x"099D4",
 50=> x"09CF6",
 51=> x"0A018",
 52=> x"0A33A",
 53=> x"0A65C",
 54=> x"0A97E",
 55=> x"0AC9F",
 56=> x"0AFC1",
 57=> x"0B2E2",
 58=> x"0B604",
 59=> x"0B925",
 60=> x"0BC46",
 61=> x"0BF67",
 62=> x"0C288",
 63=> x"0C5A9",
 64=> x"0C8C9",
 65=> x"0CBEA",
 66=> x"0CF0A",
 67=> x"0D22A",
 68=> x"0D54A",
 69=> x"0D86A",
 70=> x"0DB8A",
 71=> x"0DEAA",
 72=> x"0E1CA",
 73=> x"0E4E9",
 74=> x"0E808",
 75=> x"0EB28",
 76=> x"0EE47",
 77=> x"0F166",
 78=> x"0F484",
 79=> x"0F7A3",
 80=> x"0FAC1",
 81=> x"0FDE0",
 82=> x"100FE",
 83=> x"1041C",
 84=> x"1073A",
 85=> x"10A58",
 86=> x"10D75",
 87=> x"11092",
 88=> x"113B0",
 89=> x"116CD",
 90=> x"119EA",
 91=> x"11D06",
 92=> x"12023",
 93=> x"1233F",
 94=> x"1265B",
 95=> x"12977",
 96=> x"12C93",
 97=> x"12FAF",
 98=> x"132CA",
 99=> x"135E5",
 100=> x"13901",
 101=> x"13C1B",
 102=> x"13F36",
 103=> x"14251",
 104=> x"1456B",
 105=> x"14885",
 106=> x"14B9F",
 107=> x"14EB9",
 108=> x"151D2",
 109=> x"154EC",
 110=> x"15805",
 111=> x"15B1E",
 112=> x"15E36",
 113=> x"1614F",
 114=> x"16467",
 115=> x"1677F",
 116=> x"16A97",
 117=> x"16DAF",
 118=> x"170C6",
 119=> x"173DD",
 120=> x"176F4",
 121=> x"17A0B",
 122=> x"17D21",
 123=> x"18038",
 124=> x"1834E",
 125=> x"18664",
 126=> x"18979",
 127=> x"18C8E",
 128=> x"18FA4",
 129=> x"192B8",
 130=> x"195CD",
 131=> x"198E1",
 132=> x"19BF6",
 133=> x"19F09",
 134=> x"1A21D",
 135=> x"1A530",
 136=> x"1A844",
 137=> x"1AB56",
 138=> x"1AE69",
 139=> x"1B17B",
 140=> x"1B48D",
 141=> x"1B79F",
 142=> x"1BAB1",
 143=> x"1BDC2",
 144=> x"1C0D3",
 145=> x"1C3E4",
 146=> x"1C6F4",
 147=> x"1CA05",
 148=> x"1CD15",
 149=> x"1D024",
 150=> x"1D334",
 151=> x"1D643",
 152=> x"1D951",
 153=> x"1DC60",
 154=> x"1DF6E",
 155=> x"1E27C",
 156=> x"1E58A",
 157=> x"1E897",
 158=> x"1EBA4",
 159=> x"1EEB1",
 160=> x"1F1BD",
 161=> x"1F4CA",
 162=> x"1F7D5",
 163=> x"1FAE1",
 164=> x"1FDEC",
 165=> x"200F7",
 166=> x"20402",
 167=> x"2070C",
 168=> x"20A16",
 169=> x"20D20",
 170=> x"21029",
 171=> x"21332",
 172=> x"2163B",
 173=> x"21944",
 174=> x"21C4C",
 175=> x"21F54",
 176=> x"2225B",
 177=> x"22562",
 178=> x"22869",
 179=> x"22B6F",
 180=> x"22E75",
 181=> x"2317B",
 182=> x"23481",
 183=> x"23786",
 184=> x"23A8B",
 185=> x"23D8F",
 186=> x"24093",
 187=> x"24397",
 188=> x"2469A",
 189=> x"2499D",
 190=> x"24CA0",
 191=> x"24FA2",
 192=> x"252A4",
 193=> x"255A6",
 194=> x"258A7",
 195=> x"25BA8",
 196=> x"25EA8",
 197=> x"261A9",
 198=> x"264A8",
 199=> x"267A8",
 200=> x"26AA7",
 201=> x"26DA6",
 202=> x"270A4",
 203=> x"273A2",
 204=> x"2769F",
 205=> x"2799D",
 206=> x"27C99",
 207=> x"27F96",
 208=> x"28292",
 209=> x"2858D",
 210=> x"28889",
 211=> x"28B83",
 212=> x"28E7E",
 213=> x"29178",
 214=> x"29472",
 215=> x"2976B",
 216=> x"29A64",
 217=> x"29D5C",
 218=> x"2A054",
 219=> x"2A34C",
 220=> x"2A643",
 221=> x"2A93A",
 222=> x"2AC30",
 223=> x"2AF26",
 224=> x"2B21C",
 225=> x"2B511",
 226=> x"2B806",
 227=> x"2BAFA",
 228=> x"2BDEE",
 229=> x"2C0E2",
 230=> x"2C3D5",
 231=> x"2C6C8",
 232=> x"2C9BA",
 233=> x"2CCAC",
 234=> x"2CF9D",
 235=> x"2D28E",
 236=> x"2D57E",
 237=> x"2D86E",
 238=> x"2DB5E",
 239=> x"2DE4D",
 240=> x"2E13C",
 241=> x"2E42A",
 242=> x"2E718",
 243=> x"2EA05",
 244=> x"2ECF2",
 245=> x"2EFDF",
 246=> x"2F2CB",
 247=> x"2F5B7",
 248=> x"2F8A2",
 249=> x"2FB8C",
 250=> x"2FE77",
 251=> x"30160",
 252=> x"3044A",
 253=> x"30732",
 254=> x"30A1B",
 255=> x"30D03",
 256=> x"30FEA",
 257=> x"312D1",
 258=> x"315B8",
 259=> x"3189D",
 260=> x"31B83",
 261=> x"31E68",
 262=> x"3214D",
 263=> x"32431",
 264=> x"32714",
 265=> x"329F7",
 266=> x"32CDA",
 267=> x"32FBC",
 268=> x"3329E",
 269=> x"3357F",
 270=> x"3385F",
 271=> x"33B40",
 272=> x"33E1F",
 273=> x"340FE",
 274=> x"343DD",
 275=> x"346BB",
 276=> x"34999",
 277=> x"34C76",
 278=> x"34F53",
 279=> x"3522F",
 280=> x"3550A",
 281=> x"357E5",
 282=> x"35AC0",
 283=> x"35D9A",
 284=> x"36074",
 285=> x"3634D",
 286=> x"36625",
 287=> x"368FD",
 288=> x"36BD4",
 289=> x"36EAB",
 290=> x"37182",
 291=> x"37458",
 292=> x"3772D",
 293=> x"37A02",
 294=> x"37CD6",
 295=> x"37FAA",
 296=> x"3827D",
 297=> x"3854F",
 298=> x"38821",
 299=> x"38AF3",
 300=> x"38DC4",
 301=> x"39094",
 302=> x"39364",
 303=> x"39634",
 304=> x"39902",
 305=> x"39BD1",
 306=> x"39E9E",
 307=> x"3A16B",
 308=> x"3A438",
 309=> x"3A704",
 310=> x"3A9CF",
 311=> x"3AC9A",
 312=> x"3AF65",
 313=> x"3B22E",
 314=> x"3B4F7",
 315=> x"3B7C0",
 316=> x"3BA88",
 317=> x"3BD4F",
 318=> x"3C016",
 319=> x"3C2DD",
 320=> x"3C5A2",
 321=> x"3C867",
 322=> x"3CB2C",
 323=> x"3CDF0",
 324=> x"3D0B3",
 325=> x"3D376",
 326=> x"3D638",
 327=> x"3D8FA",
 328=> x"3DBBB",
 329=> x"3DE7B",
 330=> x"3E13B",
 331=> x"3E3FA",
 332=> x"3E6B9",
 333=> x"3E977",
 334=> x"3EC34",
 335=> x"3EEF1",
 336=> x"3F1AD",
 337=> x"3F469",
 338=> x"3F724",
 339=> x"3F9DE",
 340=> x"3FC98",
 341=> x"3FF51",
 342=> x"4020A",
 343=> x"404C1",
 344=> x"40779",
 345=> x"40A2F",
 346=> x"40CE5",
 347=> x"40F9B",
 348=> x"41250",
 349=> x"41504",
 350=> x"417B7",
 351=> x"41A6A",
 352=> x"41D1C",
 353=> x"41FCE",
 354=> x"4227F",
 355=> x"4252F",
 356=> x"427DF",
 357=> x"42A8E",
 358=> x"42D3D",
 359=> x"42FEA",
 360=> x"43298",
 361=> x"43544",
 362=> x"437F0",
 363=> x"43A9B",
 364=> x"43D46",
 365=> x"43FEF",
 366=> x"44299",
 367=> x"44541",
 368=> x"447E9",
 369=> x"44A90",
 370=> x"44D37",
 371=> x"44FDD",
 372=> x"45282",
 373=> x"45527",
 374=> x"457CB",
 375=> x"45A6E",
 376=> x"45D10",
 377=> x"45FB2",
 378=> x"46254",
 379=> x"464F4",
 380=> x"46794",
 381=> x"46A33",
 382=> x"46CD2",
 383=> x"46F70",
 384=> x"4720D",
 385=> x"474A9",
 386=> x"47745",
 387=> x"479E0",
 388=> x"47C7A",
 389=> x"47F14",
 390=> x"481AD",
 391=> x"48445",
 392=> x"486DD",
 393=> x"48974",
 394=> x"48C0A",
 395=> x"48EA0",
 396=> x"49135",
 397=> x"493C9",
 398=> x"4965C",
 399=> x"498EF",
 400=> x"49B81",
 401=> x"49E12",
 402=> x"4A0A3",
 403=> x"4A332",
 404=> x"4A5C2",
 405=> x"4A850",
 406=> x"4AADE",
 407=> x"4AD6B",
 408=> x"4AFF7",
 409=> x"4B282",
 410=> x"4B50D",
 411=> x"4B797",
 412=> x"4BA21",
 413=> x"4BCA9",
 414=> x"4BF31",
 415=> x"4C1B8",
 416=> x"4C43F",
 417=> x"4C6C5",
 418=> x"4C949",
 419=> x"4CBCE",
 420=> x"4CE51",
 421=> x"4D0D4",
 422=> x"4D356",
 423=> x"4D5D7",
 424=> x"4D858",
 425=> x"4DAD7",
 426=> x"4DD56",
 427=> x"4DFD5",
 428=> x"4E252",
 429=> x"4E4CF",
 430=> x"4E74B",
 431=> x"4E9C6",
 432=> x"4EC41",
 433=> x"4EEBA",
 434=> x"4F133",
 435=> x"4F3AB",
 436=> x"4F623",
 437=> x"4F89A",
 438=> x"4FB0F",
 439=> x"4FD85",
 440=> x"4FFF9",
 441=> x"5026D",
 442=> x"504DF",
 443=> x"50751",
 444=> x"509C3",
 445=> x"50C33",
 446=> x"50EA3",
 447=> x"51112",
 448=> x"51380",
 449=> x"515ED",
 450=> x"5185A",
 451=> x"51AC6",
 452=> x"51D31",
 453=> x"51F9B",
 454=> x"52204",
 455=> x"5246D",
 456=> x"526D5",
 457=> x"5293C",
 458=> x"52BA2",
 459=> x"52E08",
 460=> x"5306C",
 461=> x"532D0",
 462=> x"53533",
 463=> x"53795",
 464=> x"539F7",
 465=> x"53C57",
 466=> x"53EB7",
 467=> x"54116",
 468=> x"54375",
 469=> x"545D2",
 470=> x"5482F",
 471=> x"54A8A",
 472=> x"54CE5",
 473=> x"54F3F",
 474=> x"55199",
 475=> x"553F1",
 476=> x"55649",
 477=> x"558A0",
 478=> x"55AF6",
 479=> x"55D4B",
 480=> x"55F9F",
 481=> x"561F3",
 482=> x"56446",
 483=> x"56697",
 484=> x"568E8",
 485=> x"56B39",
 486=> x"56D88",
 487=> x"56FD7",
 488=> x"57224",
 489=> x"57471",
 490=> x"576BD",
 491=> x"57908",
 492=> x"57B53",
 493=> x"57D9C",
 494=> x"57FE5",
 495=> x"5822D",
 496=> x"58474",
 497=> x"586BA",
 498=> x"588FF",
 499=> x"58B43",
 500=> x"58D87",
 501=> x"58FC9",
 502=> x"5920B",
 503=> x"5944C",
 504=> x"5968C",
 505=> x"598CC",
 506=> x"59B0A",
 507=> x"59D47",
 508=> x"59F84",
 509=> x"5A1C0",
 510=> x"5A3FB",
 511=> x"5A635",
 512=> x"5A86E",
 513=> x"5AAA6",
 514=> x"5ACDE",
 515=> x"5AF14",
 516=> x"5B14A",
 517=> x"5B37E",
 518=> x"5B5B2",
 519=> x"5B7E5",
 520=> x"5BA18",
 521=> x"5BC49",
 522=> x"5BE79",
 523=> x"5C0A9",
 524=> x"5C2D7",
 525=> x"5C505",
 526=> x"5C732",
 527=> x"5C95E",
 528=> x"5CB89",
 529=> x"5CDB3",
 530=> x"5CFDC",
 531=> x"5D204",
 532=> x"5D42C",
 533=> x"5D652",
 534=> x"5D878",
 535=> x"5DA9D",
 536=> x"5DCC1",
 537=> x"5DEE4",
 538=> x"5E106",
 539=> x"5E327",
 540=> x"5E547",
 541=> x"5E766",
 542=> x"5E985",
 543=> x"5EBA2",
 544=> x"5EDBF",
 545=> x"5EFDA",
 546=> x"5F1F5",
 547=> x"5F40F",
 548=> x"5F628",
 549=> x"5F840",
 550=> x"5FA57",
 551=> x"5FC6D",
 552=> x"5FE82",
 553=> x"60096",
 554=> x"602AA",
 555=> x"604BC",
 556=> x"606CE",
 557=> x"608DE",
 558=> x"60AEE",
 559=> x"60CFD",
 560=> x"60F0A",
 561=> x"61117",
 562=> x"61323",
 563=> x"6152E",
 564=> x"61738",
 565=> x"61941",
 566=> x"61B49",
 567=> x"61D51",
 568=> x"61F57",
 569=> x"6215C",
 570=> x"62361",
 571=> x"62564",
 572=> x"62767",
 573=> x"62968",
 574=> x"62B69",
 575=> x"62D68",
 576=> x"62F67",
 577=> x"63165",
 578=> x"63361",
 579=> x"6355D",
 580=> x"63758",
 581=> x"63952",
 582=> x"63B4B",
 583=> x"63D43",
 584=> x"63F3A",
 585=> x"64130",
 586=> x"64325",
 587=> x"64519",
 588=> x"6470C",
 589=> x"648FE",
 590=> x"64AF0",
 591=> x"64CE0",
 592=> x"64ECF",
 593=> x"650BD",
 594=> x"652AB",
 595=> x"65497",
 596=> x"65683",
 597=> x"6586D",
 598=> x"65A56",
 599=> x"65C3F",
 600=> x"65E26",
 601=> x"6600D",
 602=> x"661F2",
 603=> x"663D7",
 604=> x"665BA",
 605=> x"6679D",
 606=> x"6697E",
 607=> x"66B5F",
 608=> x"66D3E",
 609=> x"66F1D",
 610=> x"670FA",
 611=> x"672D7",
 612=> x"674B3",
 613=> x"6768D",
 614=> x"67867",
 615=> x"67A3F",
 616=> x"67C17",
 617=> x"67DEE",
 618=> x"67FC3",
 619=> x"68198",
 620=> x"6836B",
 621=> x"6853E",
 622=> x"6870F",
 623=> x"688E0",
 624=> x"68AB0",
 625=> x"68C7E",
 626=> x"68E4C",
 627=> x"69018",
 628=> x"691E4",
 629=> x"693AE",
 630=> x"69578",
 631=> x"69740",
 632=> x"69908",
 633=> x"69ACE",
 634=> x"69C93",
 635=> x"69E58",
 636=> x"6A01B",
 637=> x"6A1DE",
 638=> x"6A39F",
 639=> x"6A55F",
 640=> x"6A71E",
 641=> x"6A8DD",
 642=> x"6AA9A",
 643=> x"6AC56",
 644=> x"6AE11",
 645=> x"6AFCB",
 646=> x"6B185",
 647=> x"6B33D",
 648=> x"6B4F4",
 649=> x"6B6AA",
 650=> x"6B85F",
 651=> x"6BA13",
 652=> x"6BBC5",
 653=> x"6BD77",
 654=> x"6BF28",
 655=> x"6C0D8",
 656=> x"6C287",
 657=> x"6C434",
 658=> x"6C5E1",
 659=> x"6C78D",
 660=> x"6C937",
 661=> x"6CAE1",
 662=> x"6CC89",
 663=> x"6CE30",
 664=> x"6CFD7",
 665=> x"6D17C",
 666=> x"6D320",
 667=> x"6D4C4",
 668=> x"6D666",
 669=> x"6D807",
 670=> x"6D9A7",
 671=> x"6DB46",
 672=> x"6DCE4",
 673=> x"6DE81",
 674=> x"6E01C",
 675=> x"6E1B7",
 676=> x"6E351",
 677=> x"6E4E9",
 678=> x"6E681",
 679=> x"6E817",
 680=> x"6E9AD",
 681=> x"6EB41",
 682=> x"6ECD5",
 683=> x"6EE67",
 684=> x"6EFF8",
 685=> x"6F188",
 686=> x"6F317",
 687=> x"6F4A5",
 688=> x"6F632",
 689=> x"6F7BE",
 690=> x"6F948",
 691=> x"6FAD2",
 692=> x"6FC5B",
 693=> x"6FDE2",
 694=> x"6FF68",
 695=> x"700EE",
 696=> x"70272",
 697=> x"703F5",
 698=> x"70577",
 699=> x"706F8",
 700=> x"70878",
 701=> x"709F7",
 702=> x"70B75",
 703=> x"70CF1",
 704=> x"70E6D",
 705=> x"70FE7",
 706=> x"71161",
 707=> x"712D9",
 708=> x"71450",
 709=> x"715C6",
 710=> x"7173B",
 711=> x"718AF",
 712=> x"71A22",
 713=> x"71B94",
 714=> x"71D05",
 715=> x"71E74",
 716=> x"71FE3",
 717=> x"72150",
 718=> x"722BC",
 719=> x"72427",
 720=> x"72591",
 721=> x"726FA",
 722=> x"72862",
 723=> x"729C9",
 724=> x"72B2F",
 725=> x"72C93",
 726=> x"72DF6",
 727=> x"72F59",
 728=> x"730BA",
 729=> x"7321A",
 730=> x"73379",
 731=> x"734D7",
 732=> x"73634",
 733=> x"7378F",
 734=> x"738EA",
 735=> x"73A43",
 736=> x"73B9C",
 737=> x"73CF3",
 738=> x"73E49",
 739=> x"73F9E",
 740=> x"740F2",
 741=> x"74244",
 742=> x"74396",
 743=> x"744E6",
 744=> x"74636",
 745=> x"74784",
 746=> x"748D1",
 747=> x"74A1D",
 748=> x"74B68",
 749=> x"74CB2",
 750=> x"74DFA",
 751=> x"74F42",
 752=> x"75088",
 753=> x"751CD",
 754=> x"75311",
 755=> x"75454",
 756=> x"75596",
 757=> x"756D7",
 758=> x"75816",
 759=> x"75955",
 760=> x"75A92",
 761=> x"75BCE",
 762=> x"75D09",
 763=> x"75E43",
 764=> x"75F7C",
 765=> x"760B4",
 766=> x"761EA",
 767=> x"7631F",
 768=> x"76454",
 769=> x"76587",
 770=> x"766B9",
 771=> x"767E9",
 772=> x"76919",
 773=> x"76A48",
 774=> x"76B75",
 775=> x"76CA1",
 776=> x"76DCC",
 777=> x"76EF6",
 778=> x"7701F",
 779=> x"77146",
 780=> x"7726D",
 781=> x"77392",
 782=> x"774B6",
 783=> x"775D9",
 784=> x"776FB",
 785=> x"7781C",
 786=> x"7793C",
 787=> x"77A5A",
 788=> x"77B77",
 789=> x"77C93",
 790=> x"77DAE",
 791=> x"77EC8",
 792=> x"77FE1",
 793=> x"780F8",
 794=> x"7820F",
 795=> x"78324",
 796=> x"78438",
 797=> x"7854B",
 798=> x"7865C",
 799=> x"7876D",
 800=> x"7887C",
 801=> x"7898A",
 802=> x"78A97",
 803=> x"78BA3",
 804=> x"78CAE",
 805=> x"78DB8",
 806=> x"78EC0",
 807=> x"78FC7",
 808=> x"790CD",
 809=> x"791D2",
 810=> x"792D6",
 811=> x"793D8",
 812=> x"794DA",
 813=> x"795DA",
 814=> x"796D9",
 815=> x"797D7",
 816=> x"798D4",
 817=> x"799CF",
 818=> x"79AC9",
 819=> x"79BC3",
 820=> x"79CBB",
 821=> x"79DB1",
 822=> x"79EA7",
 823=> x"79F9B",
 824=> x"7A08F",
 825=> x"7A181",
 826=> x"7A272",
 827=> x"7A362",
 828=> x"7A450",
 829=> x"7A53E",
 830=> x"7A62A",
 831=> x"7A715",
 832=> x"7A7FF",
 833=> x"7A8E7",
 834=> x"7A9CF",
 835=> x"7AAB5",
 836=> x"7AB9A",
 837=> x"7AC7E",
 838=> x"7AD61",
 839=> x"7AE43",
 840=> x"7AF23",
 841=> x"7B002",
 842=> x"7B0E0",
 843=> x"7B1BD",
 844=> x"7B299",
 845=> x"7B373",
 846=> x"7B44D",
 847=> x"7B525",
 848=> x"7B5FC",
 849=> x"7B6D1",
 850=> x"7B7A6",
 851=> x"7B879",
 852=> x"7B94B",
 853=> x"7BA1C",
 854=> x"7BAEC",
 855=> x"7BBBB",
 856=> x"7BC88",
 857=> x"7BD54",
 858=> x"7BE1F",
 859=> x"7BEE9",
 860=> x"7BFB2",
 861=> x"7C079",
 862=> x"7C13F",
 863=> x"7C204",
 864=> x"7C2C8",
 865=> x"7C38B",
 866=> x"7C44C",
 867=> x"7C50C",
 868=> x"7C5CB",
 869=> x"7C689",
 870=> x"7C746",
 871=> x"7C801",
 872=> x"7C8BB",
 873=> x"7C974",
 874=> x"7CA2C",
 875=> x"7CAE3",
 876=> x"7CB98",
 877=> x"7CC4C",
 878=> x"7CCFF",
 879=> x"7CDB1",
 880=> x"7CE62",
 881=> x"7CF11",
 882=> x"7CFBF",
 883=> x"7D06C",
 884=> x"7D118",
 885=> x"7D1C3",
 886=> x"7D26C",
 887=> x"7D314",
 888=> x"7D3BB",
 889=> x"7D461",
 890=> x"7D505",
 891=> x"7D5A9",
 892=> x"7D64B",
 893=> x"7D6EC",
 894=> x"7D78B",
 895=> x"7D82A",
 896=> x"7D8C7",
 897=> x"7D963",
 898=> x"7D9FE",
 899=> x"7DA98",
 900=> x"7DB30",
 901=> x"7DBC7",
 902=> x"7DC5E",
 903=> x"7DCF2",
 904=> x"7DD86",
 905=> x"7DE18",
 906=> x"7DEA9",
 907=> x"7DF39",
 908=> x"7DFC8",
 909=> x"7E056",
 910=> x"7E0E2",
 911=> x"7E16D",
 912=> x"7E1F7",
 913=> x"7E27F",
 914=> x"7E307",
 915=> x"7E38D",
 916=> x"7E412",
 917=> x"7E496",
 918=> x"7E518",
 919=> x"7E59A",
 920=> x"7E61A",
 921=> x"7E699",
 922=> x"7E717",
 923=> x"7E793",
 924=> x"7E80E",
 925=> x"7E888",
 926=> x"7E901",
 927=> x"7E979",
 928=> x"7E9EF",
 929=> x"7EA64",
 930=> x"7EAD8",
 931=> x"7EB4B",
 932=> x"7EBBC",
 933=> x"7EC2D",
 934=> x"7EC9C",
 935=> x"7ED09",
 936=> x"7ED76",
 937=> x"7EDE1",
 938=> x"7EE4C",
 939=> x"7EEB5",
 940=> x"7EF1C",
 941=> x"7EF83",
 942=> x"7EFE8",
 943=> x"7F04C",
 944=> x"7F0AF",
 945=> x"7F110",
 946=> x"7F171",
 947=> x"7F1D0",
 948=> x"7F22E",
 949=> x"7F28A",
 950=> x"7F2E6",
 951=> x"7F340",
 952=> x"7F399",
 953=> x"7F3F1",
 954=> x"7F447",
 955=> x"7F49D",
 956=> x"7F4F1",
 957=> x"7F544",
 958=> x"7F595",
 959=> x"7F5E6",
 960=> x"7F635",
 961=> x"7F683",
 962=> x"7F6D0",
 963=> x"7F71B",
 964=> x"7F765",
 965=> x"7F7AE",
 966=> x"7F7F6",
 967=> x"7F83D",
 968=> x"7F882",
 969=> x"7F8C6",
 970=> x"7F909",
 971=> x"7F94B",
 972=> x"7F98B",
 973=> x"7F9CA",
 974=> x"7FA08",
 975=> x"7FA45",
 976=> x"7FA80",
 977=> x"7FABB",
 978=> x"7FAF4",
 979=> x"7FB2C",
 980=> x"7FB62",
 981=> x"7FB98",
 982=> x"7FBCC",
 983=> x"7FBFF",
 984=> x"7FC30",
 985=> x"7FC61",
 986=> x"7FC90",
 987=> x"7FCBE",
 988=> x"7FCEA",
 989=> x"7FD16",
 990=> x"7FD40",
 991=> x"7FD69",
 992=> x"7FD91",
 993=> x"7FDB8",
 994=> x"7FDDD",
 995=> x"7FE01",
 996=> x"7FE24",
 997=> x"7FE45",
 998=> x"7FE66",
 999=> x"7FE85",
 1000=> x"7FEA3",
 1001=> x"7FEC0",
 1002=> x"7FEDB",
 1003=> x"7FEF5",
 1004=> x"7FF0E",
 1005=> x"7FF26",
 1006=> x"7FF3D",
 1007=> x"7FF52",
 1008=> x"7FF66",
 1009=> x"7FF79",
 1010=> x"7FF8A",
 1011=> x"7FF9B",
 1012=> x"7FFAA",
 1013=> x"7FFB8",
 1014=> x"7FFC4",
 1015=> x"7FFD0",
 1016=> x"7FFDA",
 1017=> x"7FFE3",
 1018=> x"7FFEB",
 1019=> x"7FFF1",
 1020=> x"7FFF6",
 1021=> x"7FFFA",
 1022=> x"7FFFD",
 1023=> x"7FFFF",
 1024=> x"7FFFF",
 1025=> x"7FFFE",
 1026=> x"7FFFC",
 1027=> x"7FFF8",
 1028=> x"7FFF4",
 1029=> x"7FFEE",
 1030=> x"7FFE7",
 1031=> x"7FFDF",
 1032=> x"7FFD5",
 1033=> x"7FFCA",
 1034=> x"7FFBE",
 1035=> x"7FFB1",
 1036=> x"7FFA2",
 1037=> x"7FF93",
 1038=> x"7FF82",
 1039=> x"7FF6F",
 1040=> x"7FF5C",
 1041=> x"7FF47",
 1042=> x"7FF31",
 1043=> x"7FF1A",
 1044=> x"7FF02",
 1045=> x"7FEE8",
 1046=> x"7FECE",
 1047=> x"7FEB1",
 1048=> x"7FE94",
 1049=> x"7FE76",
 1050=> x"7FE56",
 1051=> x"7FE35",
 1052=> x"7FE13",
 1053=> x"7FDEF",
 1054=> x"7FDCA",
 1055=> x"7FDA4",
 1056=> x"7FD7D",
 1057=> x"7FD55",
 1058=> x"7FD2B",
 1059=> x"7FD00",
 1060=> x"7FCD4",
 1061=> x"7FCA7",
 1062=> x"7FC78",
 1063=> x"7FC49",
 1064=> x"7FC17",
 1065=> x"7FBE5",
 1066=> x"7FBB2",
 1067=> x"7FB7D",
 1068=> x"7FB47",
 1069=> x"7FB10",
 1070=> x"7FAD7",
 1071=> x"7FA9E",
 1072=> x"7FA63",
 1073=> x"7FA27",
 1074=> x"7F9E9",
 1075=> x"7F9AB",
 1076=> x"7F96B",
 1077=> x"7F92A",
 1078=> x"7F8E8",
 1079=> x"7F8A4",
 1080=> x"7F860",
 1081=> x"7F81A",
 1082=> x"7F7D2",
 1083=> x"7F78A",
 1084=> x"7F740",
 1085=> x"7F6F5",
 1086=> x"7F6A9",
 1087=> x"7F65C",
 1088=> x"7F60D",
 1089=> x"7F5BE",
 1090=> x"7F56D",
 1091=> x"7F51A",
 1092=> x"7F4C7",
 1093=> x"7F472",
 1094=> x"7F41C",
 1095=> x"7F3C5",
 1096=> x"7F36D",
 1097=> x"7F313",
 1098=> x"7F2B8",
 1099=> x"7F25C",
 1100=> x"7F1FF",
 1101=> x"7F1A0",
 1102=> x"7F141",
 1103=> x"7F0E0",
 1104=> x"7F07E",
 1105=> x"7F01A",
 1106=> x"7EFB5",
 1107=> x"7EF50",
 1108=> x"7EEE9",
 1109=> x"7EE80",
 1110=> x"7EE17",
 1111=> x"7EDAC",
 1112=> x"7ED40",
 1113=> x"7ECD3",
 1114=> x"7EC64",
 1115=> x"7EBF5",
 1116=> x"7EB84",
 1117=> x"7EB12",
 1118=> x"7EA9E",
 1119=> x"7EA2A",
 1120=> x"7E9B4",
 1121=> x"7E93D",
 1122=> x"7E8C5",
 1123=> x"7E84B",
 1124=> x"7E7D1",
 1125=> x"7E755",
 1126=> x"7E6D8",
 1127=> x"7E65A",
 1128=> x"7E5DA",
 1129=> x"7E559",
 1130=> x"7E4D7",
 1131=> x"7E454",
 1132=> x"7E3D0",
 1133=> x"7E34A",
 1134=> x"7E2C3",
 1135=> x"7E23B",
 1136=> x"7E1B2",
 1137=> x"7E128",
 1138=> x"7E09C",
 1139=> x"7E00F",
 1140=> x"7DF81",
 1141=> x"7DEF2",
 1142=> x"7DE61",
 1143=> x"7DDCF",
 1144=> x"7DD3C",
 1145=> x"7DCA8",
 1146=> x"7DC13",
 1147=> x"7DB7C",
 1148=> x"7DAE4",
 1149=> x"7DA4B",
 1150=> x"7D9B1",
 1151=> x"7D915",
 1152=> x"7D879",
 1153=> x"7D7DB",
 1154=> x"7D73C",
 1155=> x"7D69B",
 1156=> x"7D5FA",
 1157=> x"7D557",
 1158=> x"7D4B3",
 1159=> x"7D40E",
 1160=> x"7D368",
 1161=> x"7D2C0",
 1162=> x"7D218",
 1163=> x"7D16E",
 1164=> x"7D0C2",
 1165=> x"7D016",
 1166=> x"7CF68",
 1167=> x"7CEBA",
 1168=> x"7CE0A",
 1169=> x"7CD58",
 1170=> x"7CCA6",
 1171=> x"7CBF2",
 1172=> x"7CB3E",
 1173=> x"7CA88",
 1174=> x"7C9D0",
 1175=> x"7C918",
 1176=> x"7C85E",
 1177=> x"7C7A4",
 1178=> x"7C6E8",
 1179=> x"7C62A",
 1180=> x"7C56C",
 1181=> x"7C4AC",
 1182=> x"7C3EB",
 1183=> x"7C329",
 1184=> x"7C266",
 1185=> x"7C1A2",
 1186=> x"7C0DC",
 1187=> x"7C015",
 1188=> x"7BF4D",
 1189=> x"7BE84",
 1190=> x"7BDBA",
 1191=> x"7BCEE",
 1192=> x"7BC21",
 1193=> x"7BB53",
 1194=> x"7BA84",
 1195=> x"7B9B4",
 1196=> x"7B8E2",
 1197=> x"7B810",
 1198=> x"7B73C",
 1199=> x"7B667",
 1200=> x"7B590",
 1201=> x"7B4B9",
 1202=> x"7B3E0",
 1203=> x"7B306",
 1204=> x"7B22B",
 1205=> x"7B14F",
 1206=> x"7B072",
 1207=> x"7AF93",
 1208=> x"7AEB3",
 1209=> x"7ADD2",
 1210=> x"7ACF0",
 1211=> x"7AC0D",
 1212=> x"7AB28",
 1213=> x"7AA42",
 1214=> x"7A95B",
 1215=> x"7A873",
 1216=> x"7A78A",
 1217=> x"7A6A0",
 1218=> x"7A5B4",
 1219=> x"7A4C7",
 1220=> x"7A3D9",
 1221=> x"7A2EA",
 1222=> x"7A1FA",
 1223=> x"7A108",
 1224=> x"7A015",
 1225=> x"79F21",
 1226=> x"79E2C",
 1227=> x"79D36",
 1228=> x"79C3F",
 1229=> x"79B46",
 1230=> x"79A4C",
 1231=> x"79951",
 1232=> x"79855",
 1233=> x"79758",
 1234=> x"7965A",
 1235=> x"7955A",
 1236=> x"79459",
 1237=> x"79357",
 1238=> x"79254",
 1239=> x"79150",
 1240=> x"7904A",
 1241=> x"78F44",
 1242=> x"78E3C",
 1243=> x"78D33",
 1244=> x"78C29",
 1245=> x"78B1E",
 1246=> x"78A11",
 1247=> x"78903",
 1248=> x"787F5",
 1249=> x"786E5",
 1250=> x"785D4",
 1251=> x"784C1",
 1252=> x"783AE",
 1253=> x"78299",
 1254=> x"78184",
 1255=> x"7806D",
 1256=> x"77F55",
 1257=> x"77E3B",
 1258=> x"77D21",
 1259=> x"77C06",
 1260=> x"77AE9",
 1261=> x"779CB",
 1262=> x"778AC",
 1263=> x"7778C",
 1264=> x"7766B",
 1265=> x"77548",
 1266=> x"77425",
 1267=> x"77300",
 1268=> x"771DA",
 1269=> x"770B3",
 1270=> x"76F8B",
 1271=> x"76E61",
 1272=> x"76D37",
 1273=> x"76C0B",
 1274=> x"76ADE",
 1275=> x"769B0",
 1276=> x"76881",
 1277=> x"76751",
 1278=> x"76620",
 1279=> x"764ED",
 1280=> x"763BA",
 1281=> x"76285",
 1282=> x"7614F",
 1283=> x"76018",
 1284=> x"75EE0",
 1285=> x"75DA6",
 1286=> x"75C6C",
 1287=> x"75B30",
 1288=> x"759F4",
 1289=> x"758B6",
 1290=> x"75777",
 1291=> x"75637",
 1292=> x"754F5",
 1293=> x"753B3",
 1294=> x"7526F",
 1295=> x"7512B",
 1296=> x"74FE5",
 1297=> x"74E9E",
 1298=> x"74D56",
 1299=> x"74C0D",
 1300=> x"74AC3",
 1301=> x"74977",
 1302=> x"7482B",
 1303=> x"746DD",
 1304=> x"7458E",
 1305=> x"7443E",
 1306=> x"742ED",
 1307=> x"7419B",
 1308=> x"74048",
 1309=> x"73EF3",
 1310=> x"73D9E",
 1311=> x"73C47",
 1312=> x"73AF0",
 1313=> x"73997",
 1314=> x"7383D",
 1315=> x"736E2",
 1316=> x"73585",
 1317=> x"73428",
 1318=> x"732CA",
 1319=> x"7316A",
 1320=> x"7300A",
 1321=> x"72EA8",
 1322=> x"72D45",
 1323=> x"72BE1",
 1324=> x"72A7C",
 1325=> x"72916",
 1326=> x"727AE",
 1327=> x"72646",
 1328=> x"724DD",
 1329=> x"72372",
 1330=> x"72206",
 1331=> x"72099",
 1332=> x"71F2C",
 1333=> x"71DBD",
 1334=> x"71C4C",
 1335=> x"71ADB",
 1336=> x"71969",
 1337=> x"717F6",
 1338=> x"71681",
 1339=> x"7150C",
 1340=> x"71395",
 1341=> x"7121D",
 1342=> x"710A4",
 1343=> x"70F2A",
 1344=> x"70DAF",
 1345=> x"70C33",
 1346=> x"70AB6",
 1347=> x"70938",
 1348=> x"707B8",
 1349=> x"70638",
 1350=> x"704B6",
 1351=> x"70334",
 1352=> x"701B0",
 1353=> x"7002B",
 1354=> x"6FEA5",
 1355=> x"6FD1E",
 1356=> x"6FB96",
 1357=> x"6FA0D",
 1358=> x"6F883",
 1359=> x"6F6F8",
 1360=> x"6F56C",
 1361=> x"6F3DE",
 1362=> x"6F250",
 1363=> x"6F0C0",
 1364=> x"6EF2F",
 1365=> x"6ED9E",
 1366=> x"6EC0B",
 1367=> x"6EA77",
 1368=> x"6E8E2",
 1369=> x"6E74C",
 1370=> x"6E5B5",
 1371=> x"6E41D",
 1372=> x"6E284",
 1373=> x"6E0EA",
 1374=> x"6DF4F",
 1375=> x"6DDB2",
 1376=> x"6DC15",
 1377=> x"6DA76",
 1378=> x"6D8D7",
 1379=> x"6D736",
 1380=> x"6D595",
 1381=> x"6D3F2",
 1382=> x"6D24E",
 1383=> x"6D0AA",
 1384=> x"6CF04",
 1385=> x"6CD5D",
 1386=> x"6CBB5",
 1387=> x"6CA0C",
 1388=> x"6C862",
 1389=> x"6C6B7",
 1390=> x"6C50B",
 1391=> x"6C35E",
 1392=> x"6C1AF",
 1393=> x"6C000",
 1394=> x"6BE50",
 1395=> x"6BC9E",
 1396=> x"6BAEC",
 1397=> x"6B939",
 1398=> x"6B784",
 1399=> x"6B5CF",
 1400=> x"6B418",
 1401=> x"6B261",
 1402=> x"6B0A8",
 1403=> x"6AEEE",
 1404=> x"6AD34",
 1405=> x"6AB78",
 1406=> x"6A9BB",
 1407=> x"6A7FE",
 1408=> x"6A63F",
 1409=> x"6A47F",
 1410=> x"6A2BE",
 1411=> x"6A0FC",
 1412=> x"69F3A",
 1413=> x"69D76",
 1414=> x"69BB1",
 1415=> x"699EB",
 1416=> x"69824",
 1417=> x"6965C",
 1418=> x"69493",
 1419=> x"692C9",
 1420=> x"690FE",
 1421=> x"68F32",
 1422=> x"68D65",
 1423=> x"68B97",
 1424=> x"689C8",
 1425=> x"687F8",
 1426=> x"68627",
 1427=> x"68455",
 1428=> x"68282",
 1429=> x"680AE",
 1430=> x"67ED8",
 1431=> x"67D02",
 1432=> x"67B2B",
 1433=> x"67953",
 1434=> x"6777A",
 1435=> x"675A0",
 1436=> x"673C5",
 1437=> x"671E9",
 1438=> x"6700C",
 1439=> x"66E2E",
 1440=> x"66C4F",
 1441=> x"66A6F",
 1442=> x"6688E",
 1443=> x"666AC",
 1444=> x"664C9",
 1445=> x"662E4",
 1446=> x"66100",
 1447=> x"65F1A",
 1448=> x"65D33",
 1449=> x"65B4B",
 1450=> x"65962",
 1451=> x"65778",
 1452=> x"6558D",
 1453=> x"653A1",
 1454=> x"651B4",
 1455=> x"64FC6",
 1456=> x"64DD8",
 1457=> x"64BE8",
 1458=> x"649F7",
 1459=> x"64806",
 1460=> x"64613",
 1461=> x"6441F",
 1462=> x"6422B",
 1463=> x"64035",
 1464=> x"63E3F",
 1465=> x"63C47",
 1466=> x"63A4F",
 1467=> x"63855",
 1468=> x"6365B",
 1469=> x"6345F",
 1470=> x"63263",
 1471=> x"63066",
 1472=> x"62E68",
 1473=> x"62C69",
 1474=> x"62A68",
 1475=> x"62867",
 1476=> x"62665",
 1477=> x"62462",
 1478=> x"6225F",
 1479=> x"6205A",
 1480=> x"61E54",
 1481=> x"61C4D",
 1482=> x"61A46",
 1483=> x"6183D",
 1484=> x"61633",
 1485=> x"61429",
 1486=> x"6121D",
 1487=> x"61011",
 1488=> x"60E04",
 1489=> x"60BF5",
 1490=> x"609E6",
 1491=> x"607D6",
 1492=> x"605C5",
 1493=> x"603B3",
 1494=> x"601A0",
 1495=> x"5FF8C",
 1496=> x"5FD78",
 1497=> x"5FB62",
 1498=> x"5F94B",
 1499=> x"5F734",
 1500=> x"5F51B",
 1501=> x"5F302",
 1502=> x"5F0E8",
 1503=> x"5EECD",
 1504=> x"5ECB0",
 1505=> x"5EA93",
 1506=> x"5E876",
 1507=> x"5E657",
 1508=> x"5E437",
 1509=> x"5E216",
 1510=> x"5DFF5",
 1511=> x"5DDD2",
 1512=> x"5DBAF",
 1513=> x"5D98B",
 1514=> x"5D765",
 1515=> x"5D53F",
 1516=> x"5D318",
 1517=> x"5D0F0",
 1518=> x"5CEC8",
 1519=> x"5CC9E",
 1520=> x"5CA73",
 1521=> x"5C848",
 1522=> x"5C61B",
 1523=> x"5C3EE",
 1524=> x"5C1C0",
 1525=> x"5BF91",
 1526=> x"5BD61",
 1527=> x"5BB30",
 1528=> x"5B8FF",
 1529=> x"5B6CC",
 1530=> x"5B499",
 1531=> x"5B264",
 1532=> x"5B02F",
 1533=> x"5ADF9",
 1534=> x"5ABC2",
 1535=> x"5A98A",
 1536=> x"5A751",
 1537=> x"5A518",
 1538=> x"5A2DD",
 1539=> x"5A0A2",
 1540=> x"59E66",
 1541=> x"59C29",
 1542=> x"599EB",
 1543=> x"597AC",
 1544=> x"5956C",
 1545=> x"5932C",
 1546=> x"590EA",
 1547=> x"58EA8",
 1548=> x"58C65",
 1549=> x"58A21",
 1550=> x"587DC",
 1551=> x"58597",
 1552=> x"58350",
 1553=> x"58109",
 1554=> x"57EC1",
 1555=> x"57C78",
 1556=> x"57A2E",
 1557=> x"577E3",
 1558=> x"57597",
 1559=> x"5734B",
 1560=> x"570FE",
 1561=> x"56EAF",
 1562=> x"56C60",
 1563=> x"56A11",
 1564=> x"567C0",
 1565=> x"5656F",
 1566=> x"5631C",
 1567=> x"560C9",
 1568=> x"55E75",
 1569=> x"55C20",
 1570=> x"559CB",
 1571=> x"55774",
 1572=> x"5551D",
 1573=> x"552C5",
 1574=> x"5506C",
 1575=> x"54E12",
 1576=> x"54BB8",
 1577=> x"5495D",
 1578=> x"54700",
 1579=> x"544A3",
 1580=> x"54246",
 1581=> x"53FE7",
 1582=> x"53D88",
 1583=> x"53B27",
 1584=> x"538C6",
 1585=> x"53664",
 1586=> x"53402",
 1587=> x"5319E",
 1588=> x"52F3A",
 1589=> x"52CD5",
 1590=> x"52A6F",
 1591=> x"52808",
 1592=> x"525A1",
 1593=> x"52339",
 1594=> x"520D0",
 1595=> x"51E66",
 1596=> x"51BFB",
 1597=> x"51990",
 1598=> x"51724",
 1599=> x"514B7",
 1600=> x"51249",
 1601=> x"50FDA",
 1602=> x"50D6B",
 1603=> x"50AFB",
 1604=> x"5088A",
 1605=> x"50619",
 1606=> x"503A6",
 1607=> x"50133",
 1608=> x"4FEBF",
 1609=> x"4FC4A",
 1610=> x"4F9D5",
 1611=> x"4F75E",
 1612=> x"4F4E7",
 1613=> x"4F26F",
 1614=> x"4EFF7",
 1615=> x"4ED7E",
 1616=> x"4EB03",
 1617=> x"4E889",
 1618=> x"4E60D",
 1619=> x"4E391",
 1620=> x"4E113",
 1621=> x"4DE96",
 1622=> x"4DC17",
 1623=> x"4D998",
 1624=> x"4D717",
 1625=> x"4D497",
 1626=> x"4D215",
 1627=> x"4CF93",
 1628=> x"4CD10",
 1629=> x"4CA8C",
 1630=> x"4C807",
 1631=> x"4C582",
 1632=> x"4C2FC",
 1633=> x"4C075",
 1634=> x"4BDED",
 1635=> x"4BB65",
 1636=> x"4B8DC",
 1637=> x"4B652",
 1638=> x"4B3C8",
 1639=> x"4B13D",
 1640=> x"4AEB1",
 1641=> x"4AC24",
 1642=> x"4A997",
 1643=> x"4A709",
 1644=> x"4A47A",
 1645=> x"4A1EB",
 1646=> x"49F5A",
 1647=> x"49CC9",
 1648=> x"49A38",
 1649=> x"497A6",
 1650=> x"49512",
 1651=> x"4927F",
 1652=> x"48FEA",
 1653=> x"48D55",
 1654=> x"48ABF",
 1655=> x"48829",
 1656=> x"48591",
 1657=> x"482F9",
 1658=> x"48061",
 1659=> x"47DC7",
 1660=> x"47B2D",
 1661=> x"47893",
 1662=> x"475F7",
 1663=> x"4735B",
 1664=> x"470BE",
 1665=> x"46E21",
 1666=> x"46B83",
 1667=> x"468E4",
 1668=> x"46644",
 1669=> x"463A4",
 1670=> x"46103",
 1671=> x"45E62",
 1672=> x"45BBF",
 1673=> x"4591C",
 1674=> x"45679",
 1675=> x"453D5",
 1676=> x"45130",
 1677=> x"44E8A",
 1678=> x"44BE4",
 1679=> x"4493D",
 1680=> x"44695",
 1681=> x"443ED",
 1682=> x"44144",
 1683=> x"43E9B",
 1684=> x"43BF0",
 1685=> x"43946",
 1686=> x"4369A",
 1687=> x"433EE",
 1688=> x"43141",
 1689=> x"42E94",
 1690=> x"42BE5",
 1691=> x"42937",
 1692=> x"42687",
 1693=> x"423D7",
 1694=> x"42127",
 1695=> x"41E75",
 1696=> x"41BC3",
 1697=> x"41911",
 1698=> x"4165E",
 1699=> x"413AA",
 1700=> x"410F5",
 1701=> x"40E40",
 1702=> x"40B8A",
 1703=> x"408D4",
 1704=> x"4061D",
 1705=> x"40366",
 1706=> x"400AD",
 1707=> x"3FDF5",
 1708=> x"3FB3B",
 1709=> x"3F881",
 1710=> x"3F5C6",
 1711=> x"3F30B",
 1712=> x"3F04F",
 1713=> x"3ED93",
 1714=> x"3EAD6",
 1715=> x"3E818",
 1716=> x"3E55A",
 1717=> x"3E29B",
 1718=> x"3DFDB",
 1719=> x"3DD1B",
 1720=> x"3DA5A",
 1721=> x"3D799",
 1722=> x"3D4D7",
 1723=> x"3D215",
 1724=> x"3CF52",
 1725=> x"3CC8E",
 1726=> x"3C9CA",
 1727=> x"3C705",
 1728=> x"3C440",
 1729=> x"3C17A",
 1730=> x"3BEB3",
 1731=> x"3BBEC",
 1732=> x"3B924",
 1733=> x"3B65C",
 1734=> x"3B393",
 1735=> x"3B0CA",
 1736=> x"3AE00",
 1737=> x"3AB35",
 1738=> x"3A86A",
 1739=> x"3A59E",
 1740=> x"3A2D2",
 1741=> x"3A005",
 1742=> x"39D38",
 1743=> x"39A6A",
 1744=> x"3979B",
 1745=> x"394CC",
 1746=> x"391FC",
 1747=> x"38F2C",
 1748=> x"38C5C",
 1749=> x"3898A",
 1750=> x"386B8",
 1751=> x"383E6",
 1752=> x"38113",
 1753=> x"37E40",
 1754=> x"37B6C",
 1755=> x"37897",
 1756=> x"375C2",
 1757=> x"372ED",
 1758=> x"37017",
 1759=> x"36D40",
 1760=> x"36A69",
 1761=> x"36791",
 1762=> x"364B9",
 1763=> x"361E0",
 1764=> x"35F07",
 1765=> x"35C2D",
 1766=> x"35953",
 1767=> x"35678",
 1768=> x"3539D",
 1769=> x"350C1",
 1770=> x"34DE4",
 1771=> x"34B07",
 1772=> x"3482A",
 1773=> x"3454C",
 1774=> x"3426E",
 1775=> x"33F8F",
 1776=> x"33CB0",
 1777=> x"339D0",
 1778=> x"336EF",
 1779=> x"3340E",
 1780=> x"3312D",
 1781=> x"32E4B",
 1782=> x"32B69",
 1783=> x"32886",
 1784=> x"325A3",
 1785=> x"322BF",
 1786=> x"31FDA",
 1787=> x"31CF6",
 1788=> x"31A10",
 1789=> x"3172B",
 1790=> x"31444",
 1791=> x"3115E",
 1792=> x"30E76",
 1793=> x"30B8F",
 1794=> x"308A7",
 1795=> x"305BE",
 1796=> x"302D5",
 1797=> x"2FFEC",
 1798=> x"2FD02",
 1799=> x"2FA17",
 1800=> x"2F72C",
 1801=> x"2F441",
 1802=> x"2F155",
 1803=> x"2EE69",
 1804=> x"2EB7C",
 1805=> x"2E88F",
 1806=> x"2E5A1",
 1807=> x"2E2B3",
 1808=> x"2DFC5",
 1809=> x"2DCD6",
 1810=> x"2D9E6",
 1811=> x"2D6F6",
 1812=> x"2D406",
 1813=> x"2D115",
 1814=> x"2CE24",
 1815=> x"2CB33",
 1816=> x"2C841",
 1817=> x"2C54E",
 1818=> x"2C25B",
 1819=> x"2BF68",
 1820=> x"2BC74",
 1821=> x"2B980",
 1822=> x"2B68C",
 1823=> x"2B397",
 1824=> x"2B0A1",
 1825=> x"2ADAB",
 1826=> x"2AAB5",
 1827=> x"2A7BF",
 1828=> x"2A4C8",
 1829=> x"2A1D0",
 1830=> x"29ED8",
 1831=> x"29BE0",
 1832=> x"298E7",
 1833=> x"295EE",
 1834=> x"292F5",
 1835=> x"28FFB",
 1836=> x"28D01",
 1837=> x"28A06",
 1838=> x"2870B",
 1839=> x"28410",
 1840=> x"28114",
 1841=> x"27E18",
 1842=> x"27B1B",
 1843=> x"2781E",
 1844=> x"27521",
 1845=> x"27223",
 1846=> x"26F25",
 1847=> x"26C26",
 1848=> x"26927",
 1849=> x"26628",
 1850=> x"26329",
 1851=> x"26029",
 1852=> x"25D28",
 1853=> x"25A28",
 1854=> x"25726",
 1855=> x"25425",
 1856=> x"25123",
 1857=> x"24E21",
 1858=> x"24B1F",
 1859=> x"2481C",
 1860=> x"24519",
 1861=> x"24215",
 1862=> x"23F11",
 1863=> x"23C0D",
 1864=> x"23908",
 1865=> x"23603",
 1866=> x"232FE",
 1867=> x"22FF8",
 1868=> x"22CF2",
 1869=> x"229EC",
 1870=> x"226E6",
 1871=> x"223DF",
 1872=> x"220D7",
 1873=> x"21DD0",
 1874=> x"21AC8",
 1875=> x"217BF",
 1876=> x"214B7",
 1877=> x"211AE",
 1878=> x"20EA5",
 1879=> x"20B9B",
 1880=> x"20891",
 1881=> x"20587",
 1882=> x"2027D",
 1883=> x"1FF72",
 1884=> x"1FC67",
 1885=> x"1F95B",
 1886=> x"1F650",
 1887=> x"1F344",
 1888=> x"1F037",
 1889=> x"1ED2B",
 1890=> x"1EA1E",
 1891=> x"1E710",
 1892=> x"1E403",
 1893=> x"1E0F5",
 1894=> x"1DDE7",
 1895=> x"1DAD9",
 1896=> x"1D7CA",
 1897=> x"1D4BB",
 1898=> x"1D1AC",
 1899=> x"1CE9C",
 1900=> x"1CB8D",
 1901=> x"1C87D",
 1902=> x"1C56C",
 1903=> x"1C25C",
 1904=> x"1BF4B",
 1905=> x"1BC3A",
 1906=> x"1B928",
 1907=> x"1B616",
 1908=> x"1B304",
 1909=> x"1AFF2",
 1910=> x"1ACE0",
 1911=> x"1A9CD",
 1912=> x"1A6BA",
 1913=> x"1A3A7",
 1914=> x"1A093",
 1915=> x"19D80",
 1916=> x"19A6C",
 1917=> x"19757",
 1918=> x"19443",
 1919=> x"1912E",
 1920=> x"18E19",
 1921=> x"18B04",
 1922=> x"187EE",
 1923=> x"184D9",
 1924=> x"181C3",
 1925=> x"17EAD",
 1926=> x"17B96",
 1927=> x"17880",
 1928=> x"17569",
 1929=> x"17252",
 1930=> x"16F3A",
 1931=> x"16C23",
 1932=> x"1690B",
 1933=> x"165F3",
 1934=> x"162DB",
 1935=> x"15FC3",
 1936=> x"15CAA",
 1937=> x"15991",
 1938=> x"15678",
 1939=> x"1535F",
 1940=> x"15046",
 1941=> x"14D2C",
 1942=> x"14A12",
 1943=> x"146F8",
 1944=> x"143DE",
 1945=> x"140C3",
 1946=> x"13DA9",
 1947=> x"13A8E",
 1948=> x"13773",
 1949=> x"13458",
 1950=> x"1313C",
 1951=> x"12E21",
 1952=> x"12B05",
 1953=> x"127E9",
 1954=> x"124CD",
 1955=> x"121B1",
 1956=> x"11E95",
 1957=> x"11B78",
 1958=> x"1185B",
 1959=> x"1153E",
 1960=> x"11221",
 1961=> x"10F04",
 1962=> x"10BE6",
 1963=> x"108C9",
 1964=> x"105AB",
 1965=> x"1028D",
 1966=> x"0FF6F",
 1967=> x"0FC51",
 1968=> x"0F932",
 1969=> x"0F614",
 1970=> x"0F2F5",
 1971=> x"0EFD6",
 1972=> x"0ECB7",
 1973=> x"0E998",
 1974=> x"0E679",
 1975=> x"0E359",
 1976=> x"0E03A",
 1977=> x"0DD1A",
 1978=> x"0D9FA",
 1979=> x"0D6DA",
 1980=> x"0D3BA",
 1981=> x"0D09A",
 1982=> x"0CD7A",
 1983=> x"0CA59",
 1984=> x"0C739",
 1985=> x"0C418",
 1986=> x"0C0F7",
 1987=> x"0BDD6",
 1988=> x"0BAB5",
 1989=> x"0B794",
 1990=> x"0B473",
 1991=> x"0B152",
 1992=> x"0AE30",
 1993=> x"0AB0F",
 1994=> x"0A7ED",
 1995=> x"0A4CB",
 1996=> x"0A1A9",
 1997=> x"09E87",
 1998=> x"09B65",
 1999=> x"09843",
 2000=> x"09521",
 2001=> x"091FE",
 2002=> x"08EDC",
 2003=> x"08BB9",
 2004=> x"08897",
 2005=> x"08574",
 2006=> x"08251",
 2007=> x"07F2E",
 2008=> x"07C0C",
 2009=> x"078E9",
 2010=> x"075C5",
 2011=> x"072A2",
 2012=> x"06F7F",
 2013=> x"06C5C",
 2014=> x"06938",
 2015=> x"06615",
 2016=> x"062F2",
 2017=> x"05FCE",
 2018=> x"05CAA",
 2019=> x"05987",
 2020=> x"05663",
 2021=> x"0533F",
 2022=> x"0501C",
 2023=> x"04CF8",
 2024=> x"049D4",
 2025=> x"046B0",
 2026=> x"0438C",
 2027=> x"04068",
 2028=> x"03D44",
 2029=> x"03A20",
 2030=> x"036FC",
 2031=> x"033D7",
 2032=> x"030B3",
 2033=> x"02D8F",
 2034=> x"02A6B",
 2035=> x"02746",
 2036=> x"02422",
 2037=> x"020FE",
 2038=> x"01DD9",
 2039=> x"01AB5",
 2040=> x"01791",
 2041=> x"0146C",
 2042=> x"01148",
 2043=> x"00E23",
 2044=> x"00AFF",
 2045=> x"007DB",
 2046=> x"004B6",
 2047=> x"00192",
 2048=> x"FFE6E",
 2049=> x"FFB4A",
 2050=> x"FF825",
 2051=> x"FF501",
 2052=> x"FF1DD",
 2053=> x"FEEB8",
 2054=> x"FEB94",
 2055=> x"FE86F",
 2056=> x"FE54B",
 2057=> x"FE227",
 2058=> x"FDF02",
 2059=> x"FDBDE",
 2060=> x"FD8BA",
 2061=> x"FD595",
 2062=> x"FD271",
 2063=> x"FCF4D",
 2064=> x"FCC29",
 2065=> x"FC904",
 2066=> x"FC5E0",
 2067=> x"FC2BC",
 2068=> x"FBF98",
 2069=> x"FBC74",
 2070=> x"FB950",
 2071=> x"FB62C",
 2072=> x"FB308",
 2073=> x"FAFE4",
 2074=> x"FACC1",
 2075=> x"FA99D",
 2076=> x"FA679",
 2077=> x"FA356",
 2078=> x"FA032",
 2079=> x"F9D0E",
 2080=> x"F99EB",
 2081=> x"F96C8",
 2082=> x"F93A4",
 2083=> x"F9081",
 2084=> x"F8D5E",
 2085=> x"F8A3B",
 2086=> x"F8717",
 2087=> x"F83F4",
 2088=> x"F80D2",
 2089=> x"F7DAF",
 2090=> x"F7A8C",
 2091=> x"F7769",
 2092=> x"F7447",
 2093=> x"F7124",
 2094=> x"F6E02",
 2095=> x"F6ADF",
 2096=> x"F67BD",
 2097=> x"F649B",
 2098=> x"F6179",
 2099=> x"F5E57",
 2100=> x"F5B35",
 2101=> x"F5813",
 2102=> x"F54F1",
 2103=> x"F51D0",
 2104=> x"F4EAE",
 2105=> x"F4B8D",
 2106=> x"F486C",
 2107=> x"F454B",
 2108=> x"F422A",
 2109=> x"F3F09",
 2110=> x"F3BE8",
 2111=> x"F38C7",
 2112=> x"F35A7",
 2113=> x"F3286",
 2114=> x"F2F66",
 2115=> x"F2C46",
 2116=> x"F2926",
 2117=> x"F2606",
 2118=> x"F22E6",
 2119=> x"F1FC6",
 2120=> x"F1CA7",
 2121=> x"F1987",
 2122=> x"F1668",
 2123=> x"F1349",
 2124=> x"F102A",
 2125=> x"F0D0B",
 2126=> x"F09EC",
 2127=> x"F06CE",
 2128=> x"F03AF",
 2129=> x"F0091",
 2130=> x"EFD73",
 2131=> x"EFA55",
 2132=> x"EF737",
 2133=> x"EF41A",
 2134=> x"EF0FC",
 2135=> x"EEDDF",
 2136=> x"EEAC2",
 2137=> x"EE7A5",
 2138=> x"EE488",
 2139=> x"EE16B",
 2140=> x"EDE4F",
 2141=> x"EDB33",
 2142=> x"ED817",
 2143=> x"ED4FB",
 2144=> x"ED1DF",
 2145=> x"ECEC4",
 2146=> x"ECBA8",
 2147=> x"EC88D",
 2148=> x"EC572",
 2149=> x"EC257",
 2150=> x"EBF3D",
 2151=> x"EBC22",
 2152=> x"EB908",
 2153=> x"EB5EE",
 2154=> x"EB2D4",
 2155=> x"EAFBA",
 2156=> x"EACA1",
 2157=> x"EA988",
 2158=> x"EA66F",
 2159=> x"EA356",
 2160=> x"EA03D",
 2161=> x"E9D25",
 2162=> x"E9A0D",
 2163=> x"E96F5",
 2164=> x"E93DD",
 2165=> x"E90C6",
 2166=> x"E8DAE",
 2167=> x"E8A97",
 2168=> x"E8780",
 2169=> x"E846A",
 2170=> x"E8153",
 2171=> x"E7E3D",
 2172=> x"E7B27",
 2173=> x"E7812",
 2174=> x"E74FC",
 2175=> x"E71E7",
 2176=> x"E6ED2",
 2177=> x"E6BBD",
 2178=> x"E68A9",
 2179=> x"E6594",
 2180=> x"E6280",
 2181=> x"E5F6D",
 2182=> x"E5C59",
 2183=> x"E5946",
 2184=> x"E5633",
 2185=> x"E5320",
 2186=> x"E500E",
 2187=> x"E4CFC",
 2188=> x"E49EA",
 2189=> x"E46D8",
 2190=> x"E43C6",
 2191=> x"E40B5",
 2192=> x"E3DA4",
 2193=> x"E3A94",
 2194=> x"E3783",
 2195=> x"E3473",
 2196=> x"E3164",
 2197=> x"E2E54",
 2198=> x"E2B45",
 2199=> x"E2836",
 2200=> x"E2527",
 2201=> x"E2219",
 2202=> x"E1F0B",
 2203=> x"E1BFD",
 2204=> x"E18F0",
 2205=> x"E15E2",
 2206=> x"E12D5",
 2207=> x"E0FC9",
 2208=> x"E0CBC",
 2209=> x"E09B0",
 2210=> x"E06A5",
 2211=> x"E0399",
 2212=> x"E008E",
 2213=> x"DFD83",
 2214=> x"DFA79",
 2215=> x"DF76F",
 2216=> x"DF465",
 2217=> x"DF15B",
 2218=> x"DEE52",
 2219=> x"DEB49",
 2220=> x"DE841",
 2221=> x"DE538",
 2222=> x"DE230",
 2223=> x"DDF29",
 2224=> x"DDC21",
 2225=> x"DD91A",
 2226=> x"DD614",
 2227=> x"DD30E",
 2228=> x"DD008",
 2229=> x"DCD02",
 2230=> x"DC9FD",
 2231=> x"DC6F8",
 2232=> x"DC3F3",
 2233=> x"DC0EF",
 2234=> x"DBDEB",
 2235=> x"DBAE7",
 2236=> x"DB7E4",
 2237=> x"DB4E1",
 2238=> x"DB1DF",
 2239=> x"DAEDD",
 2240=> x"DABDB",
 2241=> x"DA8DA",
 2242=> x"DA5D8",
 2243=> x"DA2D8",
 2244=> x"D9FD7",
 2245=> x"D9CD7",
 2246=> x"D99D8",
 2247=> x"D96D9",
 2248=> x"D93DA",
 2249=> x"D90DB",
 2250=> x"D8DDD",
 2251=> x"D8ADF",
 2252=> x"D87E2",
 2253=> x"D84E5",
 2254=> x"D81E8",
 2255=> x"D7EEC",
 2256=> x"D7BF0",
 2257=> x"D78F5",
 2258=> x"D75FA",
 2259=> x"D72FF",
 2260=> x"D7005",
 2261=> x"D6D0B",
 2262=> x"D6A12",
 2263=> x"D6719",
 2264=> x"D6420",
 2265=> x"D6128",
 2266=> x"D5E30",
 2267=> x"D5B38",
 2268=> x"D5841",
 2269=> x"D554B",
 2270=> x"D5255",
 2271=> x"D4F5F",
 2272=> x"D4C69",
 2273=> x"D4974",
 2274=> x"D4680",
 2275=> x"D438C",
 2276=> x"D4098",
 2277=> x"D3DA5",
 2278=> x"D3AB2",
 2279=> x"D37BF",
 2280=> x"D34CD",
 2281=> x"D31DC",
 2282=> x"D2EEB",
 2283=> x"D2BFA",
 2284=> x"D290A",
 2285=> x"D261A",
 2286=> x"D232A",
 2287=> x"D203B",
 2288=> x"D1D4D",
 2289=> x"D1A5F",
 2290=> x"D1771",
 2291=> x"D1484",
 2292=> x"D1197",
 2293=> x"D0EAB",
 2294=> x"D0BBF",
 2295=> x"D08D4",
 2296=> x"D05E9",
 2297=> x"D02FE",
 2298=> x"D0014",
 2299=> x"CFD2B",
 2300=> x"CFA42",
 2301=> x"CF759",
 2302=> x"CF471",
 2303=> x"CF18A",
 2304=> x"CEEA2",
 2305=> x"CEBBC",
 2306=> x"CE8D5",
 2307=> x"CE5F0",
 2308=> x"CE30A",
 2309=> x"CE026",
 2310=> x"CDD41",
 2311=> x"CDA5D",
 2312=> x"CD77A",
 2313=> x"CD497",
 2314=> x"CD1B5",
 2315=> x"CCED3",
 2316=> x"CCBF2",
 2317=> x"CC911",
 2318=> x"CC630",
 2319=> x"CC350",
 2320=> x"CC071",
 2321=> x"CBD92",
 2322=> x"CBAB4",
 2323=> x"CB7D6",
 2324=> x"CB4F9",
 2325=> x"CB21C",
 2326=> x"CAF3F",
 2327=> x"CAC63",
 2328=> x"CA988",
 2329=> x"CA6AD",
 2330=> x"CA3D3",
 2331=> x"CA0F9",
 2332=> x"C9E20",
 2333=> x"C9B47",
 2334=> x"C986F",
 2335=> x"C9597",
 2336=> x"C92C0",
 2337=> x"C8FE9",
 2338=> x"C8D13",
 2339=> x"C8A3E",
 2340=> x"C8769",
 2341=> x"C8494",
 2342=> x"C81C0",
 2343=> x"C7EED",
 2344=> x"C7C1A",
 2345=> x"C7948",
 2346=> x"C7676",
 2347=> x"C73A4",
 2348=> x"C70D4",
 2349=> x"C6E04",
 2350=> x"C6B34",
 2351=> x"C6865",
 2352=> x"C6596",
 2353=> x"C62C8",
 2354=> x"C5FFB",
 2355=> x"C5D2E",
 2356=> x"C5A62",
 2357=> x"C5796",
 2358=> x"C54CB",
 2359=> x"C5200",
 2360=> x"C4F36",
 2361=> x"C4C6D",
 2362=> x"C49A4",
 2363=> x"C46DC",
 2364=> x"C4414",
 2365=> x"C414D",
 2366=> x"C3E86",
 2367=> x"C3BC0",
 2368=> x"C38FB",
 2369=> x"C3636",
 2370=> x"C3372",
 2371=> x"C30AE",
 2372=> x"C2DEB",
 2373=> x"C2B29",
 2374=> x"C2867",
 2375=> x"C25A6",
 2376=> x"C22E5",
 2377=> x"C2025",
 2378=> x"C1D65",
 2379=> x"C1AA6",
 2380=> x"C17E8",
 2381=> x"C152A",
 2382=> x"C126D",
 2383=> x"C0FB1",
 2384=> x"C0CF5",
 2385=> x"C0A3A",
 2386=> x"C077F",
 2387=> x"C04C5",
 2388=> x"C020B",
 2389=> x"BFF53",
 2390=> x"BFC9A",
 2391=> x"BF9E3",
 2392=> x"BF72C",
 2393=> x"BF476",
 2394=> x"BF1C0",
 2395=> x"BEF0B",
 2396=> x"BEC56",
 2397=> x"BE9A2",
 2398=> x"BE6EF",
 2399=> x"BE43D",
 2400=> x"BE18B",
 2401=> x"BDED9",
 2402=> x"BDC29",
 2403=> x"BD979",
 2404=> x"BD6C9",
 2405=> x"BD41B",
 2406=> x"BD16C",
 2407=> x"BCEBF",
 2408=> x"BCC12",
 2409=> x"BC966",
 2410=> x"BC6BA",
 2411=> x"BC410",
 2412=> x"BC165",
 2413=> x"BBEBC",
 2414=> x"BBC13",
 2415=> x"BB96B",
 2416=> x"BB6C3",
 2417=> x"BB41C",
 2418=> x"BB176",
 2419=> x"BAED0",
 2420=> x"BAC2B",
 2421=> x"BA987",
 2422=> x"BA6E4",
 2423=> x"BA441",
 2424=> x"BA19E",
 2425=> x"B9EFD",
 2426=> x"B9C5C",
 2427=> x"B99BC",
 2428=> x"B971C",
 2429=> x"B947D",
 2430=> x"B91DF",
 2431=> x"B8F42",
 2432=> x"B8CA5",
 2433=> x"B8A09",
 2434=> x"B876D",
 2435=> x"B84D3",
 2436=> x"B8239",
 2437=> x"B7F9F",
 2438=> x"B7D07",
 2439=> x"B7A6F",
 2440=> x"B77D7",
 2441=> x"B7541",
 2442=> x"B72AB",
 2443=> x"B7016",
 2444=> x"B6D81",
 2445=> x"B6AEE",
 2446=> x"B685A",
 2447=> x"B65C8",
 2448=> x"B6337",
 2449=> x"B60A6",
 2450=> x"B5E15",
 2451=> x"B5B86",
 2452=> x"B58F7",
 2453=> x"B5669",
 2454=> x"B53DC",
 2455=> x"B514F",
 2456=> x"B4EC3",
 2457=> x"B4C38",
 2458=> x"B49AE",
 2459=> x"B4724",
 2460=> x"B449B",
 2461=> x"B4213",
 2462=> x"B3F8B",
 2463=> x"B3D04",
 2464=> x"B3A7E",
 2465=> x"B37F9",
 2466=> x"B3574",
 2467=> x"B32F0",
 2468=> x"B306D",
 2469=> x"B2DEB",
 2470=> x"B2B69",
 2471=> x"B28E9",
 2472=> x"B2668",
 2473=> x"B23E9",
 2474=> x"B216A",
 2475=> x"B1EED",
 2476=> x"B1C6F",
 2477=> x"B19F3",
 2478=> x"B1777",
 2479=> x"B14FD",
 2480=> x"B1282",
 2481=> x"B1009",
 2482=> x"B0D91",
 2483=> x"B0B19",
 2484=> x"B08A2",
 2485=> x"B062B",
 2486=> x"B03B6",
 2487=> x"B0141",
 2488=> x"AFECD",
 2489=> x"AFC5A",
 2490=> x"AF9E7",
 2491=> x"AF776",
 2492=> x"AF505",
 2493=> x"AF295",
 2494=> x"AF026",
 2495=> x"AEDB7",
 2496=> x"AEB49",
 2497=> x"AE8DC",
 2498=> x"AE670",
 2499=> x"AE405",
 2500=> x"AE19A",
 2501=> x"ADF30",
 2502=> x"ADCC7",
 2503=> x"ADA5F",
 2504=> x"AD7F8",
 2505=> x"AD591",
 2506=> x"AD32B",
 2507=> x"AD0C6",
 2508=> x"ACE62",
 2509=> x"ACBFE",
 2510=> x"AC99C",
 2511=> x"AC73A",
 2512=> x"AC4D9",
 2513=> x"AC278",
 2514=> x"AC019",
 2515=> x"ABDBA",
 2516=> x"ABB5D",
 2517=> x"AB900",
 2518=> x"AB6A3",
 2519=> x"AB448",
 2520=> x"AB1EE",
 2521=> x"AAF94",
 2522=> x"AAD3B",
 2523=> x"AAAE3",
 2524=> x"AA88C",
 2525=> x"AA635",
 2526=> x"AA3E0",
 2527=> x"AA18B",
 2528=> x"A9F37",
 2529=> x"A9CE4",
 2530=> x"A9A91",
 2531=> x"A9840",
 2532=> x"A95EF",
 2533=> x"A93A0",
 2534=> x"A9151",
 2535=> x"A8F02",
 2536=> x"A8CB5",
 2537=> x"A8A69",
 2538=> x"A881D",
 2539=> x"A85D2",
 2540=> x"A8388",
 2541=> x"A813F",
 2542=> x"A7EF7",
 2543=> x"A7CB0",
 2544=> x"A7A69",
 2545=> x"A7824",
 2546=> x"A75DF",
 2547=> x"A739B",
 2548=> x"A7158",
 2549=> x"A6F16",
 2550=> x"A6CD4",
 2551=> x"A6A94",
 2552=> x"A6854",
 2553=> x"A6615",
 2554=> x"A63D7",
 2555=> x"A619A",
 2556=> x"A5F5E",
 2557=> x"A5D23",
 2558=> x"A5AE8",
 2559=> x"A58AF",
 2560=> x"A5676",
 2561=> x"A543E",
 2562=> x"A5207",
 2563=> x"A4FD1",
 2564=> x"A4D9C",
 2565=> x"A4B67",
 2566=> x"A4934",
 2567=> x"A4701",
 2568=> x"A44D0",
 2569=> x"A429F",
 2570=> x"A406F",
 2571=> x"A3E40",
 2572=> x"A3C12",
 2573=> x"A39E5",
 2574=> x"A37B8",
 2575=> x"A358D",
 2576=> x"A3362",
 2577=> x"A3138",
 2578=> x"A2F10",
 2579=> x"A2CE8",
 2580=> x"A2AC1",
 2581=> x"A289B",
 2582=> x"A2675",
 2583=> x"A2451",
 2584=> x"A222E",
 2585=> x"A200B",
 2586=> x"A1DEA",
 2587=> x"A1BC9",
 2588=> x"A19A9",
 2589=> x"A178A",
 2590=> x"A156D",
 2591=> x"A1350",
 2592=> x"A1133",
 2593=> x"A0F18",
 2594=> x"A0CFE",
 2595=> x"A0AE5",
 2596=> x"A08CC",
 2597=> x"A06B5",
 2598=> x"A049E",
 2599=> x"A0288",
 2600=> x"A0074",
 2601=> x"9FE60",
 2602=> x"9FC4D",
 2603=> x"9FA3B",
 2604=> x"9F82A",
 2605=> x"9F61A",
 2606=> x"9F40B",
 2607=> x"9F1FC",
 2608=> x"9EFEF",
 2609=> x"9EDE3",
 2610=> x"9EBD7",
 2611=> x"9E9CD",
 2612=> x"9E7C3",
 2613=> x"9E5BA",
 2614=> x"9E3B3",
 2615=> x"9E1AC",
 2616=> x"9DFA6",
 2617=> x"9DDA1",
 2618=> x"9DB9E",
 2619=> x"9D99B",
 2620=> x"9D799",
 2621=> x"9D598",
 2622=> x"9D397",
 2623=> x"9D198",
 2624=> x"9CF9A",
 2625=> x"9CD9D",
 2626=> x"9CBA1",
 2627=> x"9C9A5",
 2628=> x"9C7AB",
 2629=> x"9C5B1",
 2630=> x"9C3B9",
 2631=> x"9C1C1",
 2632=> x"9BFCB",
 2633=> x"9BDD5",
 2634=> x"9BBE1",
 2635=> x"9B9ED",
 2636=> x"9B7FA",
 2637=> x"9B609",
 2638=> x"9B418",
 2639=> x"9B228",
 2640=> x"9B03A",
 2641=> x"9AE4C",
 2642=> x"9AC5F",
 2643=> x"9AA73",
 2644=> x"9A888",
 2645=> x"9A69E",
 2646=> x"9A4B5",
 2647=> x"9A2CD",
 2648=> x"9A0E6",
 2649=> x"99F00",
 2650=> x"99D1C",
 2651=> x"99B37",
 2652=> x"99954",
 2653=> x"99772",
 2654=> x"99591",
 2655=> x"993B1",
 2656=> x"991D2",
 2657=> x"98FF4",
 2658=> x"98E17",
 2659=> x"98C3B",
 2660=> x"98A60",
 2661=> x"98886",
 2662=> x"986AD",
 2663=> x"984D5",
 2664=> x"982FE",
 2665=> x"98128",
 2666=> x"97F52",
 2667=> x"97D7E",
 2668=> x"97BAB",
 2669=> x"979D9",
 2670=> x"97808",
 2671=> x"97638",
 2672=> x"97469",
 2673=> x"9729B",
 2674=> x"970CE",
 2675=> x"96F02",
 2676=> x"96D37",
 2677=> x"96B6D",
 2678=> x"969A4",
 2679=> x"967DC",
 2680=> x"96615",
 2681=> x"9644F",
 2682=> x"9628A",
 2683=> x"960C6",
 2684=> x"95F04",
 2685=> x"95D42",
 2686=> x"95B81",
 2687=> x"959C1",
 2688=> x"95802",
 2689=> x"95645",
 2690=> x"95488",
 2691=> x"952CC",
 2692=> x"95112",
 2693=> x"94F58",
 2694=> x"94D9F",
 2695=> x"94BE8",
 2696=> x"94A31",
 2697=> x"9487C",
 2698=> x"946C7",
 2699=> x"94514",
 2700=> x"94362",
 2701=> x"941B0",
 2702=> x"94000",
 2703=> x"93E51",
 2704=> x"93CA2",
 2705=> x"93AF5",
 2706=> x"93949",
 2707=> x"9379E",
 2708=> x"935F4",
 2709=> x"9344B",
 2710=> x"932A3",
 2711=> x"930FC",
 2712=> x"92F56",
 2713=> x"92DB2",
 2714=> x"92C0E",
 2715=> x"92A6B",
 2716=> x"928CA",
 2717=> x"92729",
 2718=> x"9258A",
 2719=> x"923EB",
 2720=> x"9224E",
 2721=> x"920B1",
 2722=> x"91F16",
 2723=> x"91D7C",
 2724=> x"91BE3",
 2725=> x"91A4B",
 2726=> x"918B4",
 2727=> x"9171E",
 2728=> x"91589",
 2729=> x"913F5",
 2730=> x"91262",
 2731=> x"910D1",
 2732=> x"90F40",
 2733=> x"90DB0",
 2734=> x"90C22",
 2735=> x"90A94",
 2736=> x"90908",
 2737=> x"9077D",
 2738=> x"905F3",
 2739=> x"9046A",
 2740=> x"902E2",
 2741=> x"9015B",
 2742=> x"8FFD5",
 2743=> x"8FE50",
 2744=> x"8FCCC",
 2745=> x"8FB4A",
 2746=> x"8F9C8",
 2747=> x"8F848",
 2748=> x"8F6C8",
 2749=> x"8F54A",
 2750=> x"8F3CD",
 2751=> x"8F251",
 2752=> x"8F0D6",
 2753=> x"8EF5C",
 2754=> x"8EDE3",
 2755=> x"8EC6B",
 2756=> x"8EAF4",
 2757=> x"8E97F",
 2758=> x"8E80A",
 2759=> x"8E697",
 2760=> x"8E525",
 2761=> x"8E3B4",
 2762=> x"8E243",
 2763=> x"8E0D4",
 2764=> x"8DF67",
 2765=> x"8DDFA",
 2766=> x"8DC8E",
 2767=> x"8DB23",
 2768=> x"8D9BA",
 2769=> x"8D852",
 2770=> x"8D6EA",
 2771=> x"8D584",
 2772=> x"8D41F",
 2773=> x"8D2BB",
 2774=> x"8D158",
 2775=> x"8CFF6",
 2776=> x"8CE96",
 2777=> x"8CD36",
 2778=> x"8CBD8",
 2779=> x"8CA7B",
 2780=> x"8C91E",
 2781=> x"8C7C3",
 2782=> x"8C669",
 2783=> x"8C510",
 2784=> x"8C3B9",
 2785=> x"8C262",
 2786=> x"8C10D",
 2787=> x"8BFB8",
 2788=> x"8BE65",
 2789=> x"8BD13",
 2790=> x"8BBC2",
 2791=> x"8BA72",
 2792=> x"8B923",
 2793=> x"8B7D5",
 2794=> x"8B689",
 2795=> x"8B53D",
 2796=> x"8B3F3",
 2797=> x"8B2AA",
 2798=> x"8B162",
 2799=> x"8B01B",
 2800=> x"8AED5",
 2801=> x"8AD91",
 2802=> x"8AC4D",
 2803=> x"8AB0B",
 2804=> x"8A9C9",
 2805=> x"8A889",
 2806=> x"8A74A",
 2807=> x"8A60C",
 2808=> x"8A4D0",
 2809=> x"8A394",
 2810=> x"8A25A",
 2811=> x"8A120",
 2812=> x"89FE8",
 2813=> x"89EB1",
 2814=> x"89D7B",
 2815=> x"89C46",
 2816=> x"89B13",
 2817=> x"899E0",
 2818=> x"898AF",
 2819=> x"8977F",
 2820=> x"89650",
 2821=> x"89522",
 2822=> x"893F5",
 2823=> x"892C9",
 2824=> x"8919F",
 2825=> x"89075",
 2826=> x"88F4D",
 2827=> x"88E26",
 2828=> x"88D00",
 2829=> x"88BDB",
 2830=> x"88AB8",
 2831=> x"88995",
 2832=> x"88874",
 2833=> x"88754",
 2834=> x"88635",
 2835=> x"88517",
 2836=> x"883FA",
 2837=> x"882DF",
 2838=> x"881C5",
 2839=> x"880AB",
 2840=> x"87F93",
 2841=> x"87E7C",
 2842=> x"87D67",
 2843=> x"87C52",
 2844=> x"87B3F",
 2845=> x"87A2C",
 2846=> x"8791B",
 2847=> x"8780B",
 2848=> x"876FD",
 2849=> x"875EF",
 2850=> x"874E2",
 2851=> x"873D7",
 2852=> x"872CD",
 2853=> x"871C4",
 2854=> x"870BC",
 2855=> x"86FB6",
 2856=> x"86EB0",
 2857=> x"86DAC",
 2858=> x"86CA9",
 2859=> x"86BA7",
 2860=> x"86AA6",
 2861=> x"869A6",
 2862=> x"868A8",
 2863=> x"867AB",
 2864=> x"866AF",
 2865=> x"865B4",
 2866=> x"864BA",
 2867=> x"863C1",
 2868=> x"862CA",
 2869=> x"861D4",
 2870=> x"860DF",
 2871=> x"85FEB",
 2872=> x"85EF8",
 2873=> x"85E06",
 2874=> x"85D16",
 2875=> x"85C27",
 2876=> x"85B39",
 2877=> x"85A4C",
 2878=> x"85960",
 2879=> x"85876",
 2880=> x"8578D",
 2881=> x"856A5",
 2882=> x"855BE",
 2883=> x"854D8",
 2884=> x"853F3",
 2885=> x"85310",
 2886=> x"8522E",
 2887=> x"8514D",
 2888=> x"8506D",
 2889=> x"84F8E",
 2890=> x"84EB1",
 2891=> x"84DD5",
 2892=> x"84CFA",
 2893=> x"84C20",
 2894=> x"84B47",
 2895=> x"84A70",
 2896=> x"84999",
 2897=> x"848C4",
 2898=> x"847F0",
 2899=> x"8471E",
 2900=> x"8464C",
 2901=> x"8457C",
 2902=> x"844AD",
 2903=> x"843DF",
 2904=> x"84312",
 2905=> x"84246",
 2906=> x"8417C",
 2907=> x"840B3",
 2908=> x"83FEB",
 2909=> x"83F24",
 2910=> x"83E5E",
 2911=> x"83D9A",
 2912=> x"83CD7",
 2913=> x"83C15",
 2914=> x"83B54",
 2915=> x"83A94",
 2916=> x"839D6",
 2917=> x"83918",
 2918=> x"8385C",
 2919=> x"837A2",
 2920=> x"836E8",
 2921=> x"83630",
 2922=> x"83578",
 2923=> x"834C2",
 2924=> x"8340E",
 2925=> x"8335A",
 2926=> x"832A8",
 2927=> x"831F6",
 2928=> x"83146",
 2929=> x"83098",
 2930=> x"82FEA",
 2931=> x"82F3E",
 2932=> x"82E92",
 2933=> x"82DE8",
 2934=> x"82D40",
 2935=> x"82C98",
 2936=> x"82BF2",
 2937=> x"82B4D",
 2938=> x"82AA9",
 2939=> x"82A06",
 2940=> x"82965",
 2941=> x"828C4",
 2942=> x"82825",
 2943=> x"82787",
 2944=> x"826EB",
 2945=> x"8264F",
 2946=> x"825B5",
 2947=> x"8251C",
 2948=> x"82484",
 2949=> x"823ED",
 2950=> x"82358",
 2951=> x"822C4",
 2952=> x"82231",
 2953=> x"8219F",
 2954=> x"8210E",
 2955=> x"8207F",
 2956=> x"81FF1",
 2957=> x"81F64",
 2958=> x"81ED8",
 2959=> x"81E4E",
 2960=> x"81DC5",
 2961=> x"81D3D",
 2962=> x"81CB6",
 2963=> x"81C30",
 2964=> x"81BAC",
 2965=> x"81B29",
 2966=> x"81AA7",
 2967=> x"81A26",
 2968=> x"819A6",
 2969=> x"81928",
 2970=> x"818AB",
 2971=> x"8182F",
 2972=> x"817B5",
 2973=> x"8173B",
 2974=> x"816C3",
 2975=> x"8164C",
 2976=> x"815D6",
 2977=> x"81562",
 2978=> x"814EE",
 2979=> x"8147C",
 2980=> x"8140B",
 2981=> x"8139C",
 2982=> x"8132D",
 2983=> x"812C0",
 2984=> x"81254",
 2985=> x"811E9",
 2986=> x"81180",
 2987=> x"81117",
 2988=> x"810B0",
 2989=> x"8104B",
 2990=> x"80FE6",
 2991=> x"80F82",
 2992=> x"80F20",
 2993=> x"80EBF",
 2994=> x"80E60",
 2995=> x"80E01",
 2996=> x"80DA4",
 2997=> x"80D48",
 2998=> x"80CED",
 2999=> x"80C93",
 3000=> x"80C3B",
 3001=> x"80BE4",
 3002=> x"80B8E",
 3003=> x"80B39",
 3004=> x"80AE6",
 3005=> x"80A93",
 3006=> x"80A42",
 3007=> x"809F3",
 3008=> x"809A4",
 3009=> x"80957",
 3010=> x"8090B",
 3011=> x"808C0",
 3012=> x"80876",
 3013=> x"8082E",
 3014=> x"807E6",
 3015=> x"807A0",
 3016=> x"8075C",
 3017=> x"80718",
 3018=> x"806D6",
 3019=> x"80695",
 3020=> x"80655",
 3021=> x"80617",
 3022=> x"805D9",
 3023=> x"8059D",
 3024=> x"80562",
 3025=> x"80529",
 3026=> x"804F0",
 3027=> x"804B9",
 3028=> x"80483",
 3029=> x"8044E",
 3030=> x"8041B",
 3031=> x"803E9",
 3032=> x"803B7",
 3033=> x"80388",
 3034=> x"80359",
 3035=> x"8032C",
 3036=> x"80300",
 3037=> x"802D5",
 3038=> x"802AB",
 3039=> x"80283",
 3040=> x"8025C",
 3041=> x"80236",
 3042=> x"80211",
 3043=> x"801ED",
 3044=> x"801CB",
 3045=> x"801AA",
 3046=> x"8018A",
 3047=> x"8016C",
 3048=> x"8014F",
 3049=> x"80132",
 3050=> x"80118",
 3051=> x"800FE",
 3052=> x"800E6",
 3053=> x"800CF",
 3054=> x"800B9",
 3055=> x"800A4",
 3056=> x"80091",
 3057=> x"8007E",
 3058=> x"8006D",
 3059=> x"8005E",
 3060=> x"8004F",
 3061=> x"80042",
 3062=> x"80036",
 3063=> x"8002B",
 3064=> x"80021",
 3065=> x"80019",
 3066=> x"80012",
 3067=> x"8000C",
 3068=> x"80008",
 3069=> x"80004",
 3070=> x"80002",
 3071=> x"80001",
 3072=> x"80001",
 3073=> x"80003",
 3074=> x"80006",
 3075=> x"8000A",
 3076=> x"8000F",
 3077=> x"80015",
 3078=> x"8001D",
 3079=> x"80026",
 3080=> x"80030",
 3081=> x"8003C",
 3082=> x"80048",
 3083=> x"80056",
 3084=> x"80065",
 3085=> x"80076",
 3086=> x"80087",
 3087=> x"8009A",
 3088=> x"800AE",
 3089=> x"800C3",
 3090=> x"800DA",
 3091=> x"800F2",
 3092=> x"8010B",
 3093=> x"80125",
 3094=> x"80140",
 3095=> x"8015D",
 3096=> x"8017B",
 3097=> x"8019A",
 3098=> x"801BB",
 3099=> x"801DC",
 3100=> x"801FF",
 3101=> x"80223",
 3102=> x"80248",
 3103=> x"8026F",
 3104=> x"80297",
 3105=> x"802C0",
 3106=> x"802EA",
 3107=> x"80316",
 3108=> x"80342",
 3109=> x"80370",
 3110=> x"8039F",
 3111=> x"803D0",
 3112=> x"80401",
 3113=> x"80434",
 3114=> x"80468",
 3115=> x"8049E",
 3116=> x"804D4",
 3117=> x"8050C",
 3118=> x"80545",
 3119=> x"80580",
 3120=> x"805BB",
 3121=> x"805F8",
 3122=> x"80636",
 3123=> x"80675",
 3124=> x"806B5",
 3125=> x"806F7",
 3126=> x"8073A",
 3127=> x"8077E",
 3128=> x"807C3",
 3129=> x"8080A",
 3130=> x"80852",
 3131=> x"8089B",
 3132=> x"808E5",
 3133=> x"80930",
 3134=> x"8097D",
 3135=> x"809CB",
 3136=> x"80A1A",
 3137=> x"80A6B",
 3138=> x"80ABC",
 3139=> x"80B0F",
 3140=> x"80B63",
 3141=> x"80BB9",
 3142=> x"80C0F",
 3143=> x"80C67",
 3144=> x"80CC0",
 3145=> x"80D1A",
 3146=> x"80D76",
 3147=> x"80DD2",
 3148=> x"80E30",
 3149=> x"80E8F",
 3150=> x"80EF0",
 3151=> x"80F51",
 3152=> x"80FB4",
 3153=> x"81018",
 3154=> x"8107D",
 3155=> x"810E4",
 3156=> x"8114B",
 3157=> x"811B4",
 3158=> x"8121F",
 3159=> x"8128A",
 3160=> x"812F7",
 3161=> x"81364",
 3162=> x"813D3",
 3163=> x"81444",
 3164=> x"814B5",
 3165=> x"81528",
 3166=> x"8159C",
 3167=> x"81611",
 3168=> x"81687",
 3169=> x"816FF",
 3170=> x"81778",
 3171=> x"817F2",
 3172=> x"8186D",
 3173=> x"818E9",
 3174=> x"81967",
 3175=> x"819E6",
 3176=> x"81A66",
 3177=> x"81AE8",
 3178=> x"81B6A",
 3179=> x"81BEE",
 3180=> x"81C73",
 3181=> x"81CF9",
 3182=> x"81D81",
 3183=> x"81E09",
 3184=> x"81E93",
 3185=> x"81F1E",
 3186=> x"81FAA",
 3187=> x"82038",
 3188=> x"820C7",
 3189=> x"82157",
 3190=> x"821E8",
 3191=> x"8227A",
 3192=> x"8230E",
 3193=> x"823A2",
 3194=> x"82439",
 3195=> x"824D0",
 3196=> x"82568",
 3197=> x"82602",
 3198=> x"8269D",
 3199=> x"82739",
 3200=> x"827D6",
 3201=> x"82875",
 3202=> x"82914",
 3203=> x"829B5",
 3204=> x"82A57",
 3205=> x"82AFB",
 3206=> x"82B9F",
 3207=> x"82C45",
 3208=> x"82CEC",
 3209=> x"82D94",
 3210=> x"82E3D",
 3211=> x"82EE8",
 3212=> x"82F94",
 3213=> x"83041",
 3214=> x"830EF",
 3215=> x"8319E",
 3216=> x"8324F",
 3217=> x"83301",
 3218=> x"833B4",
 3219=> x"83468",
 3220=> x"8351D",
 3221=> x"835D4",
 3222=> x"8368C",
 3223=> x"83745",
 3224=> x"837FF",
 3225=> x"838BA",
 3226=> x"83977",
 3227=> x"83A35",
 3228=> x"83AF4",
 3229=> x"83BB4",
 3230=> x"83C75",
 3231=> x"83D38",
 3232=> x"83DFC",
 3233=> x"83EC1",
 3234=> x"83F87",
 3235=> x"8404E",
 3236=> x"84117",
 3237=> x"841E1",
 3238=> x"842AC",
 3239=> x"84378",
 3240=> x"84445",
 3241=> x"84514",
 3242=> x"845E4",
 3243=> x"846B5",
 3244=> x"84787",
 3245=> x"8485A",
 3246=> x"8492F",
 3247=> x"84A04",
 3248=> x"84ADB",
 3249=> x"84BB3",
 3250=> x"84C8D",
 3251=> x"84D67",
 3252=> x"84E43",
 3253=> x"84F20",
 3254=> x"84FFE",
 3255=> x"850DD",
 3256=> x"851BD",
 3257=> x"8529F",
 3258=> x"85382",
 3259=> x"85466",
 3260=> x"8554B",
 3261=> x"85631",
 3262=> x"85719",
 3263=> x"85801",
 3264=> x"858EB",
 3265=> x"859D6",
 3266=> x"85AC2",
 3267=> x"85BB0",
 3268=> x"85C9E",
 3269=> x"85D8E",
 3270=> x"85E7F",
 3271=> x"85F71",
 3272=> x"86065",
 3273=> x"86159",
 3274=> x"8624F",
 3275=> x"86345",
 3276=> x"8643D",
 3277=> x"86537",
 3278=> x"86631",
 3279=> x"8672C",
 3280=> x"86829",
 3281=> x"86927",
 3282=> x"86A26",
 3283=> x"86B26",
 3284=> x"86C28",
 3285=> x"86D2A",
 3286=> x"86E2E",
 3287=> x"86F33",
 3288=> x"87039",
 3289=> x"87140",
 3290=> x"87248",
 3291=> x"87352",
 3292=> x"8745D",
 3293=> x"87569",
 3294=> x"87676",
 3295=> x"87784",
 3296=> x"87893",
 3297=> x"879A4",
 3298=> x"87AB5",
 3299=> x"87BC8",
 3300=> x"87CDC",
 3301=> x"87DF1",
 3302=> x"87F08",
 3303=> x"8801F",
 3304=> x"88138",
 3305=> x"88252",
 3306=> x"8836D",
 3307=> x"88489",
 3308=> x"885A6",
 3309=> x"886C4",
 3310=> x"887E4",
 3311=> x"88905",
 3312=> x"88A27",
 3313=> x"88B4A",
 3314=> x"88C6E",
 3315=> x"88D93",
 3316=> x"88EBA",
 3317=> x"88FE1",
 3318=> x"8910A",
 3319=> x"89234",
 3320=> x"8935F",
 3321=> x"8948B",
 3322=> x"895B8",
 3323=> x"896E7",
 3324=> x"89817",
 3325=> x"89947",
 3326=> x"89A79",
 3327=> x"89BAC",
 3328=> x"89CE1",
 3329=> x"89E16",
 3330=> x"89F4C",
 3331=> x"8A084",
 3332=> x"8A1BD",
 3333=> x"8A2F7",
 3334=> x"8A432",
 3335=> x"8A56E",
 3336=> x"8A6AB",
 3337=> x"8A7EA",
 3338=> x"8A929",
 3339=> x"8AA6A",
 3340=> x"8ABAC",
 3341=> x"8ACEF",
 3342=> x"8AE33",
 3343=> x"8AF78",
 3344=> x"8B0BE",
 3345=> x"8B206",
 3346=> x"8B34E",
 3347=> x"8B498",
 3348=> x"8B5E3",
 3349=> x"8B72F",
 3350=> x"8B87C",
 3351=> x"8B9CA",
 3352=> x"8BB1A",
 3353=> x"8BC6A",
 3354=> x"8BDBC",
 3355=> x"8BF0E",
 3356=> x"8C062",
 3357=> x"8C1B7",
 3358=> x"8C30D",
 3359=> x"8C464",
 3360=> x"8C5BD",
 3361=> x"8C716",
 3362=> x"8C871",
 3363=> x"8C9CC",
 3364=> x"8CB29",
 3365=> x"8CC87",
 3366=> x"8CDE6",
 3367=> x"8CF46",
 3368=> x"8D0A7",
 3369=> x"8D20A",
 3370=> x"8D36D",
 3371=> x"8D4D1",
 3372=> x"8D637",
 3373=> x"8D79E",
 3374=> x"8D906",
 3375=> x"8DA6F",
 3376=> x"8DBD9",
 3377=> x"8DD44",
 3378=> x"8DEB0",
 3379=> x"8E01D",
 3380=> x"8E18C",
 3381=> x"8E2FB",
 3382=> x"8E46C",
 3383=> x"8E5DE",
 3384=> x"8E751",
 3385=> x"8E8C5",
 3386=> x"8EA3A",
 3387=> x"8EBB0",
 3388=> x"8ED27",
 3389=> x"8EE9F",
 3390=> x"8F019",
 3391=> x"8F193",
 3392=> x"8F30F",
 3393=> x"8F48B",
 3394=> x"8F609",
 3395=> x"8F788",
 3396=> x"8F908",
 3397=> x"8FA89",
 3398=> x"8FC0B",
 3399=> x"8FD8E",
 3400=> x"8FF12",
 3401=> x"90098",
 3402=> x"9021E",
 3403=> x"903A5",
 3404=> x"9052E",
 3405=> x"906B8",
 3406=> x"90842",
 3407=> x"909CE",
 3408=> x"90B5B",
 3409=> x"90CE9",
 3410=> x"90E78",
 3411=> x"91008",
 3412=> x"91199",
 3413=> x"9132B",
 3414=> x"914BF",
 3415=> x"91653",
 3416=> x"917E9",
 3417=> x"9197F",
 3418=> x"91B17",
 3419=> x"91CAF",
 3420=> x"91E49",
 3421=> x"91FE4",
 3422=> x"9217F",
 3423=> x"9231C",
 3424=> x"924BA",
 3425=> x"92659",
 3426=> x"927F9",
 3427=> x"9299A",
 3428=> x"92B3C",
 3429=> x"92CE0",
 3430=> x"92E84",
 3431=> x"93029",
 3432=> x"931D0",
 3433=> x"93377",
 3434=> x"9351F",
 3435=> x"936C9",
 3436=> x"93873",
 3437=> x"93A1F",
 3438=> x"93BCC",
 3439=> x"93D79",
 3440=> x"93F28",
 3441=> x"940D8",
 3442=> x"94289",
 3443=> x"9443B",
 3444=> x"945ED",
 3445=> x"947A1",
 3446=> x"94956",
 3447=> x"94B0C",
 3448=> x"94CC3",
 3449=> x"94E7B",
 3450=> x"95035",
 3451=> x"951EF",
 3452=> x"953AA",
 3453=> x"95566",
 3454=> x"95723",
 3455=> x"958E2",
 3456=> x"95AA1",
 3457=> x"95C61",
 3458=> x"95E22",
 3459=> x"95FE5",
 3460=> x"961A8",
 3461=> x"9636D",
 3462=> x"96532",
 3463=> x"966F8",
 3464=> x"968C0",
 3465=> x"96A88",
 3466=> x"96C52",
 3467=> x"96E1C",
 3468=> x"96FE8",
 3469=> x"971B4",
 3470=> x"97382",
 3471=> x"97550",
 3472=> x"97720",
 3473=> x"978F1",
 3474=> x"97AC2",
 3475=> x"97C95",
 3476=> x"97E68",
 3477=> x"9803D",
 3478=> x"98212",
 3479=> x"983E9",
 3480=> x"985C1",
 3481=> x"98799",
 3482=> x"98973",
 3483=> x"98B4D",
 3484=> x"98D29",
 3485=> x"98F06",
 3486=> x"990E3",
 3487=> x"992C2",
 3488=> x"994A1",
 3489=> x"99682",
 3490=> x"99863",
 3491=> x"99A46",
 3492=> x"99C29",
 3493=> x"99E0E",
 3494=> x"99FF3",
 3495=> x"9A1DA",
 3496=> x"9A3C1",
 3497=> x"9A5AA",
 3498=> x"9A793",
 3499=> x"9A97D",
 3500=> x"9AB69",
 3501=> x"9AD55",
 3502=> x"9AF43",
 3503=> x"9B131",
 3504=> x"9B320",
 3505=> x"9B510",
 3506=> x"9B702",
 3507=> x"9B8F4",
 3508=> x"9BAE7",
 3509=> x"9BCDB",
 3510=> x"9BED0",
 3511=> x"9C0C6",
 3512=> x"9C2BD",
 3513=> x"9C4B5",
 3514=> x"9C6AE",
 3515=> x"9C8A8",
 3516=> x"9CAA3",
 3517=> x"9CC9F",
 3518=> x"9CE9B",
 3519=> x"9D099",
 3520=> x"9D298",
 3521=> x"9D497",
 3522=> x"9D698",
 3523=> x"9D899",
 3524=> x"9DA9C",
 3525=> x"9DC9F",
 3526=> x"9DEA4",
 3527=> x"9E0A9",
 3528=> x"9E2AF",
 3529=> x"9E4B7",
 3530=> x"9E6BF",
 3531=> x"9E8C8",
 3532=> x"9EAD2",
 3533=> x"9ECDD",
 3534=> x"9EEE9",
 3535=> x"9F0F6",
 3536=> x"9F303",
 3537=> x"9F512",
 3538=> x"9F722",
 3539=> x"9F932",
 3540=> x"9FB44",
 3541=> x"9FD56",
 3542=> x"9FF6A",
 3543=> x"A017E",
 3544=> x"A0393",
 3545=> x"A05A9",
 3546=> x"A07C0",
 3547=> x"A09D8",
 3548=> x"A0BF1",
 3549=> x"A0E0B",
 3550=> x"A1026",
 3551=> x"A1241",
 3552=> x"A145E",
 3553=> x"A167B",
 3554=> x"A189A",
 3555=> x"A1AB9",
 3556=> x"A1CD9",
 3557=> x"A1EFA",
 3558=> x"A211C",
 3559=> x"A233F",
 3560=> x"A2563",
 3561=> x"A2788",
 3562=> x"A29AE",
 3563=> x"A2BD4",
 3564=> x"A2DFC",
 3565=> x"A3024",
 3566=> x"A324D",
 3567=> x"A3477",
 3568=> x"A36A2",
 3569=> x"A38CE",
 3570=> x"A3AFB",
 3571=> x"A3D29",
 3572=> x"A3F57",
 3573=> x"A4187",
 3574=> x"A43B7",
 3575=> x"A45E8",
 3576=> x"A481B",
 3577=> x"A4A4E",
 3578=> x"A4C82",
 3579=> x"A4EB6",
 3580=> x"A50EC",
 3581=> x"A5322",
 3582=> x"A555A",
 3583=> x"A5792",
 3584=> x"A59CB",
 3585=> x"A5C05",
 3586=> x"A5E40",
 3587=> x"A607C",
 3588=> x"A62B9",
 3589=> x"A64F6",
 3590=> x"A6734",
 3591=> x"A6974",
 3592=> x"A6BB4",
 3593=> x"A6DF5",
 3594=> x"A7037",
 3595=> x"A7279",
 3596=> x"A74BD",
 3597=> x"A7701",
 3598=> x"A7946",
 3599=> x"A7B8C",
 3600=> x"A7DD3",
 3601=> x"A801B",
 3602=> x"A8264",
 3603=> x"A84AD",
 3604=> x"A86F8",
 3605=> x"A8943",
 3606=> x"A8B8F",
 3607=> x"A8DDC",
 3608=> x"A9029",
 3609=> x"A9278",
 3610=> x"A94C7",
 3611=> x"A9718",
 3612=> x"A9969",
 3613=> x"A9BBA",
 3614=> x"A9E0D",
 3615=> x"AA061",
 3616=> x"AA2B5",
 3617=> x"AA50A",
 3618=> x"AA760",
 3619=> x"AA9B7",
 3620=> x"AAC0F",
 3621=> x"AAE67",
 3622=> x"AB0C1",
 3623=> x"AB31B",
 3624=> x"AB576",
 3625=> x"AB7D1",
 3626=> x"ABA2E",
 3627=> x"ABC8B",
 3628=> x"ABEEA",
 3629=> x"AC149",
 3630=> x"AC3A9",
 3631=> x"AC609",
 3632=> x"AC86B",
 3633=> x"ACACD",
 3634=> x"ACD30",
 3635=> x"ACF94",
 3636=> x"AD1F8",
 3637=> x"AD45E",
 3638=> x"AD6C4",
 3639=> x"AD92B",
 3640=> x"ADB93",
 3641=> x"ADDFC",
 3642=> x"AE065",
 3643=> x"AE2CF",
 3644=> x"AE53A",
 3645=> x"AE7A6",
 3646=> x"AEA13",
 3647=> x"AEC80",
 3648=> x"AEEEE",
 3649=> x"AF15D",
 3650=> x"AF3CD",
 3651=> x"AF63D",
 3652=> x"AF8AF",
 3653=> x"AFB21",
 3654=> x"AFD93",
 3655=> x"B0007",
 3656=> x"B027B",
 3657=> x"B04F1",
 3658=> x"B0766",
 3659=> x"B09DD",
 3660=> x"B0C55",
 3661=> x"B0ECD",
 3662=> x"B1146",
 3663=> x"B13BF",
 3664=> x"B163A",
 3665=> x"B18B5",
 3666=> x"B1B31",
 3667=> x"B1DAE",
 3668=> x"B202B",
 3669=> x"B22AA",
 3670=> x"B2529",
 3671=> x"B27A8",
 3672=> x"B2A29",
 3673=> x"B2CAA",
 3674=> x"B2F2C",
 3675=> x"B31AF",
 3676=> x"B3432",
 3677=> x"B36B7",
 3678=> x"B393B",
 3679=> x"B3BC1",
 3680=> x"B3E48",
 3681=> x"B40CF",
 3682=> x"B4357",
 3683=> x"B45DF",
 3684=> x"B4869",
 3685=> x"B4AF3",
 3686=> x"B4D7E",
 3687=> x"B5009",
 3688=> x"B5295",
 3689=> x"B5522",
 3690=> x"B57B0",
 3691=> x"B5A3E",
 3692=> x"B5CCE",
 3693=> x"B5F5D",
 3694=> x"B61EE",
 3695=> x"B647F",
 3696=> x"B6711",
 3697=> x"B69A4",
 3698=> x"B6C37",
 3699=> x"B6ECB",
 3700=> x"B7160",
 3701=> x"B73F6",
 3702=> x"B768C",
 3703=> x"B7923",
 3704=> x"B7BBB",
 3705=> x"B7E53",
 3706=> x"B80EC",
 3707=> x"B8386",
 3708=> x"B8620",
 3709=> x"B88BB",
 3710=> x"B8B57",
 3711=> x"B8DF3",
 3712=> x"B9090",
 3713=> x"B932E",
 3714=> x"B95CD",
 3715=> x"B986C",
 3716=> x"B9B0C",
 3717=> x"B9DAC",
 3718=> x"BA04E",
 3719=> x"BA2F0",
 3720=> x"BA592",
 3721=> x"BA835",
 3722=> x"BAAD9",
 3723=> x"BAD7E",
 3724=> x"BB023",
 3725=> x"BB2C9",
 3726=> x"BB570",
 3727=> x"BB817",
 3728=> x"BBABF",
 3729=> x"BBD67",
 3730=> x"BC011",
 3731=> x"BC2BA",
 3732=> x"BC565",
 3733=> x"BC810",
 3734=> x"BCABC",
 3735=> x"BCD68",
 3736=> x"BD016",
 3737=> x"BD2C3",
 3738=> x"BD572",
 3739=> x"BD821",
 3740=> x"BDAD1",
 3741=> x"BDD81",
 3742=> x"BE032",
 3743=> x"BE2E4",
 3744=> x"BE596",
 3745=> x"BE849",
 3746=> x"BEAFC",
 3747=> x"BEDB0",
 3748=> x"BF065",
 3749=> x"BF31B",
 3750=> x"BF5D1",
 3751=> x"BF887",
 3752=> x"BFB3F",
 3753=> x"BFDF6",
 3754=> x"C00AF",
 3755=> x"C0368",
 3756=> x"C0622",
 3757=> x"C08DC",
 3758=> x"C0B97",
 3759=> x"C0E53",
 3760=> x"C110F",
 3761=> x"C13CC",
 3762=> x"C1689",
 3763=> x"C1947",
 3764=> x"C1C06",
 3765=> x"C1EC5",
 3766=> x"C2185",
 3767=> x"C2445",
 3768=> x"C2706",
 3769=> x"C29C8",
 3770=> x"C2C8A",
 3771=> x"C2F4D",
 3772=> x"C3210",
 3773=> x"C34D4",
 3774=> x"C3799",
 3775=> x"C3A5E",
 3776=> x"C3D23",
 3777=> x"C3FEA",
 3778=> x"C42B1",
 3779=> x"C4578",
 3780=> x"C4840",
 3781=> x"C4B09",
 3782=> x"C4DD2",
 3783=> x"C509B",
 3784=> x"C5366",
 3785=> x"C5631",
 3786=> x"C58FC",
 3787=> x"C5BC8",
 3788=> x"C5E95",
 3789=> x"C6162",
 3790=> x"C642F",
 3791=> x"C66FE",
 3792=> x"C69CC",
 3793=> x"C6C9C",
 3794=> x"C6F6C",
 3795=> x"C723C",
 3796=> x"C750D",
 3797=> x"C77DF",
 3798=> x"C7AB1",
 3799=> x"C7D83",
 3800=> x"C8056",
 3801=> x"C832A",
 3802=> x"C85FE",
 3803=> x"C88D3",
 3804=> x"C8BA8",
 3805=> x"C8E7E",
 3806=> x"C9155",
 3807=> x"C942C",
 3808=> x"C9703",
 3809=> x"C99DB",
 3810=> x"C9CB3",
 3811=> x"C9F8C",
 3812=> x"CA266",
 3813=> x"CA540",
 3814=> x"CA81B",
 3815=> x"CAAF6",
 3816=> x"CADD1",
 3817=> x"CB0AD",
 3818=> x"CB38A",
 3819=> x"CB667",
 3820=> x"CB945",
 3821=> x"CBC23",
 3822=> x"CBF02",
 3823=> x"CC1E1",
 3824=> x"CC4C0",
 3825=> x"CC7A1",
 3826=> x"CCA81",
 3827=> x"CCD62",
 3828=> x"CD044",
 3829=> x"CD326",
 3830=> x"CD609",
 3831=> x"CD8EC",
 3832=> x"CDBCF",
 3833=> x"CDEB3",
 3834=> x"CE198",
 3835=> x"CE47D",
 3836=> x"CE763",
 3837=> x"CEA48",
 3838=> x"CED2F",
 3839=> x"CF016",
 3840=> x"CF2FD",
 3841=> x"CF5E5",
 3842=> x"CF8CE",
 3843=> x"CFBB6",
 3844=> x"CFEA0",
 3845=> x"D0189",
 3846=> x"D0474",
 3847=> x"D075E",
 3848=> x"D0A49",
 3849=> x"D0D35",
 3850=> x"D1021",
 3851=> x"D130E",
 3852=> x"D15FB",
 3853=> x"D18E8",
 3854=> x"D1BD6",
 3855=> x"D1EC4",
 3856=> x"D21B3",
 3857=> x"D24A2",
 3858=> x"D2792",
 3859=> x"D2A82",
 3860=> x"D2D72",
 3861=> x"D3063",
 3862=> x"D3354",
 3863=> x"D3646",
 3864=> x"D3938",
 3865=> x"D3C2B",
 3866=> x"D3F1E",
 3867=> x"D4212",
 3868=> x"D4506",
 3869=> x"D47FA",
 3870=> x"D4AEF",
 3871=> x"D4DE4",
 3872=> x"D50DA",
 3873=> x"D53D0",
 3874=> x"D56C6",
 3875=> x"D59BD",
 3876=> x"D5CB4",
 3877=> x"D5FAC",
 3878=> x"D62A4",
 3879=> x"D659C",
 3880=> x"D6895",
 3881=> x"D6B8E",
 3882=> x"D6E88",
 3883=> x"D7182",
 3884=> x"D747D",
 3885=> x"D7777",
 3886=> x"D7A73",
 3887=> x"D7D6E",
 3888=> x"D806A",
 3889=> x"D8367",
 3890=> x"D8663",
 3891=> x"D8961",
 3892=> x"D8C5E",
 3893=> x"D8F5C",
 3894=> x"D925A",
 3895=> x"D9559",
 3896=> x"D9858",
 3897=> x"D9B58",
 3898=> x"D9E57",
 3899=> x"DA158",
 3900=> x"DA458",
 3901=> x"DA759",
 3902=> x"DAA5A",
 3903=> x"DAD5C",
 3904=> x"DB05E",
 3905=> x"DB360",
 3906=> x"DB663",
 3907=> x"DB966",
 3908=> x"DBC69",
 3909=> x"DBF6D",
 3910=> x"DC271",
 3911=> x"DC575",
 3912=> x"DC87A",
 3913=> x"DCB7F",
 3914=> x"DCE85",
 3915=> x"DD18B",
 3916=> x"DD491",
 3917=> x"DD797",
 3918=> x"DDA9E",
 3919=> x"DDDA5",
 3920=> x"DE0AC",
 3921=> x"DE3B4",
 3922=> x"DE6BC",
 3923=> x"DE9C5",
 3924=> x"DECCE",
 3925=> x"DEFD7",
 3926=> x"DF2E0",
 3927=> x"DF5EA",
 3928=> x"DF8F4",
 3929=> x"DFBFE",
 3930=> x"DFF09",
 3931=> x"E0214",
 3932=> x"E051F",
 3933=> x"E082B",
 3934=> x"E0B36",
 3935=> x"E0E43",
 3936=> x"E114F",
 3937=> x"E145C",
 3938=> x"E1769",
 3939=> x"E1A76",
 3940=> x"E1D84",
 3941=> x"E2092",
 3942=> x"E23A0",
 3943=> x"E26AF",
 3944=> x"E29BD",
 3945=> x"E2CCC",
 3946=> x"E2FDC",
 3947=> x"E32EB",
 3948=> x"E35FB",
 3949=> x"E390C",
 3950=> x"E3C1C",
 3951=> x"E3F2D",
 3952=> x"E423E",
 3953=> x"E454F",
 3954=> x"E4861",
 3955=> x"E4B73",
 3956=> x"E4E85",
 3957=> x"E5197",
 3958=> x"E54AA",
 3959=> x"E57BC",
 3960=> x"E5AD0",
 3961=> x"E5DE3",
 3962=> x"E60F7",
 3963=> x"E640A",
 3964=> x"E671F",
 3965=> x"E6A33",
 3966=> x"E6D48",
 3967=> x"E705C",
 3968=> x"E7372",
 3969=> x"E7687",
 3970=> x"E799C",
 3971=> x"E7CB2",
 3972=> x"E7FC8",
 3973=> x"E82DF",
 3974=> x"E85F5",
 3975=> x"E890C",
 3976=> x"E8C23",
 3977=> x"E8F3A",
 3978=> x"E9251",
 3979=> x"E9569",
 3980=> x"E9881",
 3981=> x"E9B99",
 3982=> x"E9EB1",
 3983=> x"EA1CA",
 3984=> x"EA4E2",
 3985=> x"EA7FB",
 3986=> x"EAB14",
 3987=> x"EAE2E",
 3988=> x"EB147",
 3989=> x"EB461",
 3990=> x"EB77B",
 3991=> x"EBA95",
 3992=> x"EBDAF",
 3993=> x"EC0CA",
 3994=> x"EC3E5",
 3995=> x"EC6FF",
 3996=> x"ECA1B",
 3997=> x"ECD36",
 3998=> x"ED051",
 3999=> x"ED36D",
 4000=> x"ED689",
 4001=> x"ED9A5",
 4002=> x"EDCC1",
 4003=> x"EDFDD",
 4004=> x"EE2FA",
 4005=> x"EE616",
 4006=> x"EE933",
 4007=> x"EEC50",
 4008=> x"EEF6E",
 4009=> x"EF28B",
 4010=> x"EF5A8",
 4011=> x"EF8C6",
 4012=> x"EFBE4",
 4013=> x"EFF02",
 4014=> x"F0220",
 4015=> x"F053F",
 4016=> x"F085D",
 4017=> x"F0B7C",
 4018=> x"F0E9A",
 4019=> x"F11B9",
 4020=> x"F14D8",
 4021=> x"F17F8",
 4022=> x"F1B17",
 4023=> x"F1E36",
 4024=> x"F2156",
 4025=> x"F2476",
 4026=> x"F2796",
 4027=> x"F2AB6",
 4028=> x"F2DD6",
 4029=> x"F30F6",
 4030=> x"F3416",
 4031=> x"F3737",
 4032=> x"F3A57",
 4033=> x"F3D78",
 4034=> x"F4099",
 4035=> x"F43BA",
 4036=> x"F46DB",
 4037=> x"F49FC",
 4038=> x"F4D1E",
 4039=> x"F503F",
 4040=> x"F5361",
 4041=> x"F5682",
 4042=> x"F59A4",
 4043=> x"F5CC6",
 4044=> x"F5FE8",
 4045=> x"F630A",
 4046=> x"F662C",
 4047=> x"F694E",
 4048=> x"F6C70",
 4049=> x"F6F93",
 4050=> x"F72B5",
 4051=> x"F75D8",
 4052=> x"F78FB",
 4053=> x"F7C1D",
 4054=> x"F7F40",
 4055=> x"F8263",
 4056=> x"F8586",
 4057=> x"F88A9",
 4058=> x"F8BCC",
 4059=> x"F8EEF",
 4060=> x"F9213",
 4061=> x"F9536",
 4062=> x"F9859",
 4063=> x"F9B7D",
 4064=> x"F9EA0",
 4065=> x"FA1C4",
 4066=> x"FA4E7",
 4067=> x"FA80B",
 4068=> x"FAB2F",
 4069=> x"FAE53",
 4070=> x"FB176",
 4071=> x"FB49A",
 4072=> x"FB7BE",
 4073=> x"FBAE2",
 4074=> x"FBE06",
 4075=> x"FC12A",
 4076=> x"FC44E",
 4077=> x"FC772",
 4078=> x"FCA97",
 4079=> x"FCDBB",
 4080=> x"FD0DF",
 4081=> x"FD403",
 4082=> x"FD727",
 4083=> x"FDA4C",
 4084=> x"FDD70",
 4085=> x"FE094",
 4086=> x"FE3B9",
 4087=> x"FE6DD",
 4088=> x"FEA02",
 4089=> x"FED26",
 4090=> x"FF04A",
 4091=> x"FF36F",
 4092=> x"FF693",
 4093=> x"FF9B8",
 4094=> x"FFCDC",
 4095=> x"00000");

begin

process (clk)
begin-- process
if clk'event and clk = '1' then
DOUT_aux<=memoria(to_integer(unsigned(addr)));
end if;
end process;
DOUT<=DOUT_aux(19 downto 2)&"00";
end rtl;
