
library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity decoder_epp is
  port (
    CLK : in  std_logic;c_vector (1 downto 0));
end;

architecture rtl of decoder_epp is

begin


end rtl;
